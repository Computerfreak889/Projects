PK
     ąnY�|oy[ y[    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23":["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2"],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27":["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3"],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29":[],"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-neg":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-pos":[],"pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-neg":[],"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23"],"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1":["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21"],"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2":["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19"],"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27"],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0":["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13"],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1":["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12"],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23"],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27"],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_4":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_5":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_6":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_7":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_8":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_9":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_10":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_11":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_12":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_13":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_14":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_15":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_16":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_17":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_18":[],"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_19":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_0":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_1":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_2":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_3":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23"],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_5":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27"],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_7":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_8":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_9":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_10":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_11":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12":["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1"],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13":["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0"],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_14":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_15":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_16":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_17":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_18":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19":["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2"],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_20":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21":["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1"],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_22":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_23":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_24":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_25":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_26":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_27":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_28":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_29":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_30":[],"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_31":[]},"pin_to_color":{"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23":"#FF937E","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27":"#001544","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29":"#000000","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-neg":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-pos":"#000000","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-neg":"#000000","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0":"#FF937E","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1":"#005F39","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2":"#95003A","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3":"#001544","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0":"#010067","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1":"#9E008E","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2":"#FF937E","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3":"#001544","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_4":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_5":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_6":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_7":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_8":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_9":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_10":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_11":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_12":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_13":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_14":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_15":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_16":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_17":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_18":"#000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_19":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_0":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_1":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_2":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_3":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4":"#FF937E","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_5":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6":"#001544","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_7":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_8":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_9":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_10":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_11":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12":"#9E008E","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13":"#010067","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_14":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_15":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_16":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_17":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_18":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19":"#95003A","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_20":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21":"#005F39","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_22":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_23":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_24":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_25":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_26":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_27":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_28":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_29":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_30":"#000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_31":"#000000"},"pin_to_state":{"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29":"neutral","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-neg":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-pos":"neutral","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-neg":"neutral","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0":"neutral","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1":"neutral","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2":"neutral","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_4":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_5":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_6":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_7":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_8":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_9":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_10":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_11":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_12":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_13":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_14":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_15":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_16":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_17":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_18":"neutral","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_19":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_0":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_1":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_2":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_3":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_5":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_7":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_8":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_9":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_10":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_11":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_14":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_15":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_16":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_17":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_18":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_20":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_22":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_23":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_24":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_25":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_26":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_27":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_28":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_29":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_30":"neutral","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_31":"neutral"},"next_color_idx":8,"wires_placed_in_order":[["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13"],["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12"],["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4"],["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6"],["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21"],["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19"],["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23"],["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0"],["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2"],["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27"],["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3"],["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13"]]],[[],[["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12"]]],[[],[["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4"]]],[[],[["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6"]]],[[],[["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21"]]],[[],[["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19"]]],[[["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2"]],[]],[[],[["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23"]]],[[],[["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0"]]],[[],[["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2"]]],[[["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3"]],[]],[[],[["pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27"]]],[[],[["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3"]]],[[],[["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23":"0000000000000002","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27":"0000000000000003","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29":"_","pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_0_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_0_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_1_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_1_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_2_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_2_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_3_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_3_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_4_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_4_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_5_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_5_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_6_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_6_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_7_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_7_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_8_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_8_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_9_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_9_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_10_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_10_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_11_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_11_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_12_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_12_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_13_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_13_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_14_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_14_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_15_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_15_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_16_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_16_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_17_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_17_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_18_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_18_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_19_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_19_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_20_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_20_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_21_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_21_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_22_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_22_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_23_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_24_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_24_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_25_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_25_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_26_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_26_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_27_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_28_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_28_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_0_29_polarity-neg":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-pos":"_","pin-type-power-rail_309183b8-21a3-4c1e-b571-ced0cd74321a_1_29_polarity-neg":"_","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0":"0000000000000002","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1":"0000000000000004","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2":"0000000000000005","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3":"0000000000000003","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0":"0000000000000000","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1":"0000000000000001","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2":"0000000000000002","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3":"0000000000000003","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_4":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_5":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_6":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_7":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_8":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_9":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_10":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_11":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_12":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_13":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_14":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_15":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_16":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_17":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_18":"_","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_19":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_0":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_1":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_2":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_3":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4":"0000000000000002","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_5":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6":"0000000000000003","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_7":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_8":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_9":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_10":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_11":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12":"0000000000000001","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13":"0000000000000000","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_14":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_15":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_16":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_17":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_18":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19":"0000000000000005","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_20":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21":"0000000000000004","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_22":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_23":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_24":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_25":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_26":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_27":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_28":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_29":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_30":"_","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_31":"_"},"component_id_to_pins":{"c7b3b410-08ac-4775-976d-255d687d29f7":["0","1","2","3"],"8900e024-6b2c-4d26-a66e-08abec8766f9":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19"],"6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13"],"0000000000000001":["pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12"],"0000000000000004":["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21"],"0000000000000005":["pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19"],"0000000000000002":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2"],"0000000000000003":["pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27","pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6","pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3","pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000002":"Net 2","0000000000000003":"Net 3"},"all_breadboard_info_list":["2eae479a-c502-4024-b039-df95f0384e84_63_2_True_205_-170.00000000000003_up","309183b8-21a3-4c1e-b571-ced0cd74321a_30_2_True_535_220_up"],"breadboard_info_list":["309183b8-21a3-4c1e-b571-ced0cd74321a_30_2_True_535_220_up"],"componentsData":[{"compProperties":{},"position":[595.4916625000001,14.067411499999992],"typeId":"d38bde87-c312-441a-8093-b1322deb823a","componentVersion":1,"instanceId":"c7b3b410-08ac-4775-976d-255d687d29f7","orientation":"up","circleData":[[572.5,65.00000000000001],[587.4319090000001,65.41474099999995],[602.3638195000001,64.585199],[618.5400205000001,65.41474699999993]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[81.25,402.5],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7","orientation":"up","circleData":[[62.5,545],[77.5,545],[92.5,545],[107.5,545],[122.50000000000017,545],[137.50000000000017,545],[152.50000000000017,545],[167.50000000000017,545],[197.50000000000017,545],[212.5000000000001,545],[227.5000000000001,545],[242.5000000000001,545],[257.5000000000001,545],[272.5000000000001,545],[8.5,260],[23.499999999999886,260],[38.5,260],[53.5,260],[68.5,260],[83.5,260],[98.5,260],[113.5000000000001,260],[128.50000000000017,260],[143.5000000000001,260],[167.50000000000017,260],[182.5000000000001,260],[197.50000000000017,260],[212.5000000000001,260],[227.5000000000001,260],[242.5000000000001,260],[257.5000000000001,260],[272.5000000000001,260]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"98363baf-1e93-495d-bc05-59cfbf1a3583\",\"explorerHtmlId\":\"5080dacc-1b7d-4353-b02d-6d54b6516599\",\"nameHtmlId\":\"e8a8de26-dc3a-4764-9173-223c3587553d\",\"nameInputHtmlId\":\"46100c8f-e217-457f-8b58-8e9ec7ff5ef6\",\"explorerChildHtmlId\":\"78e01b94-3763-4cab-9a50-bc39e982bd39\",\"explorerCarrotOpenHtmlId\":\"f384916b-af2e-4527-8984-81fbf697b2f6\",\"explorerCarrotClosedHtmlId\":\"958d0d47-b2f5-4b1c-a5a0-614b3eb674f3\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"1225fffc-d7b5-4987-b165-46ff4f53c3ed\",\"explorerHtmlId\":\"27b7b099-b287-4cb2-8d69-de1b59e6bfce\",\"nameHtmlId\":\"82b1b6de-7335-49f7-9ef3-cc760adefbaf\",\"nameInputHtmlId\":\"8faae78b-b28c-4954-a70d-9cfee045b989\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"34b6c8b4-96b1-4f6f-b1b9-6cdf7b698cf2\",\"explorerHtmlId\":\"a78017ba-640e-43f8-9f01-49c32e088618\",\"nameHtmlId\":\"6f3811da-bede-4f75-88ae-9d2fe38f52ed\",\"nameInputHtmlId\":\"1f690d9d-c919-4f22-b945-2d3625e8b0b2\",\"code\":\"\"},0,","codeLabelPosition":[81.25000000000001,245.00000000000006],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[32.25625299999987,5.837631500000043],"typeId":"12011600-a4b1-4790-940a-709c15856539","componentVersion":1,"instanceId":"8900e024-6b2c-4d26-a66e-08abec8766f9","orientation":"down","circleData":[[272.5,35.00000000000001],[272.5,50.00000000000002],[272.5,65],[272.5,79.99999999999997],[227.50000000000006,102.49999999999997],[212.50000000000006,102.49999999999997],[197.50000000000006,102.49999999999997],[182.49999999999983,102.49999999999997],[167.49999999999983,102.49999999999997],[152.49999999999983,102.50000000000003],[137.49999999999986,102.49999999999997],[122.49999999999986,102.49999999999997],[107.49999999999986,102.49999999999997],[92.49999999999989,102.49999999999997],[77.49999999999989,102.49999999999997],[62.499999999999886,102.49999999999997],[47.499999999999915,102.49999999999997],[32.49999999999993,102.49999999999991],[17.499999999999922,102.49999999999991],[2.499999999999922,102.49999999999991]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-110.46159","left":"-213.96420","width":"955.28266","height":"782.96159","x":"-213.96420","y":"-110.46159"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13\",\"endPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0\",\"rawStartPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_13\",\"rawEndPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"272.5000000000_545.0000000000\\\",\\\"272.5000000000_590.0000000000\\\",\\\"332.5000000000_590.0000000000\\\",\\\"332.5000000000_35.0000000000\\\",\\\"272.5000000000_35.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12\",\"endPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1\",\"rawStartPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_12\",\"rawEndPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"257.5000000000_545.0000000000\\\",\\\"257.5000000000_605.0000000000\\\",\\\"347.5000000000_605.0000000000\\\",\\\"347.5000000000_50.0000000000\\\",\\\"272.5000000000_50.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21\",\"endPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1\",\"rawStartPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_21\",\"rawEndPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"113.5000000000_260.0000000000\\\",\\\"113.5000000000_241.2500000000\\\",\\\"115.0000000000_241.2500000000\\\",\\\"115.0000000000_170.0000000000\\\",\\\"542.5000000000_170.0000000000\\\",\\\"542.5000000000_110.2073705000\\\",\\\"587.4319090000_110.2073705000\\\",\\\"587.4319090000_65.4147410000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19\",\"endPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2\",\"rawStartPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_19\",\"rawEndPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"83.5000000000_260.0000000000\\\",\\\"83.5000000000_241.2500000000\\\",\\\"85.0000000000_241.2500000000\\\",\\\"85.0000000000_177.5000000000\\\",\\\"557.5000000000_177.5000000000\\\",\\\"557.5000000000_109.7925995000\\\",\\\"602.3638195000_109.7925995000\\\",\\\"602.3638195000_64.5851990000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23\",\"endPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_0\",\"rawEndPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"497.5000000000_575.0000000000\\\",\\\"497.5000000000_620.0000000000\\\",\\\"122.5000000000_620.0000000000\\\",\\\"122.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23\",\"endPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_2\",\"rawEndPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"527.5000000000_575.0000000000\\\",\\\"527.5000000000_140.0000000000\\\",\\\"377.5000000000_140.0000000000\\\",\\\"377.5000000000_65.0000000000\\\",\\\"272.5000000000_65.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23\",\"endPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_309183b8-21a3-4c1e-b571-ced0cd74321a_0_23_1\",\"rawEndPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"512.5000000000_575.0000000000\\\",\\\"512.5000000000_125.0000000000\\\",\\\"572.5000000000_125.0000000000\\\",\\\"572.5000000000_65.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27\",\"endPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_0\",\"rawEndPinId\":\"pin-type-component_6c1f6bf3-7f94-4f9f-8d33-5eddd381a9d7_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"497.5000000000_635.0000000000\\\",\\\"152.5000000000_635.0000000000\\\",\\\"152.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27\",\"endPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_1\",\"rawEndPinId\":\"pin-type-component_8900e024-6b2c-4d26-a66e-08abec8766f9_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"512.5000000000_635.0000000000\\\",\\\"512.5000000000_590.0000000000\\\",\\\"392.5000000000_590.0000000000\\\",\\\"392.5000000000_80.0000000000\\\",\\\"272.5000000000_80.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-breadboard_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27\",\"endPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_309183b8-21a3-4c1e-b571-ced0cd74321a_0_27_2\",\"rawEndPinId\":\"pin-type-component_c7b3b410-08ac-4775-976d-255d687d29f7_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"527.5000000000_635.0000000000\\\",\\\"572.5000000000_635.0000000000\\\",\\\"572.5000000000_110.2073735000\\\",\\\"618.5400205000_110.2073735000\\\",\\\"618.5400205000_65.4147470000\\\"]}\"}"],"projectDescription":""}PK
     ąnY               jsons/PK
     ąnYc�E�  �     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Ultrasonic Sensor","category":["User Defined"],"id":"d38bde87-c312-441a-8093-b1322deb823a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c49e1bc-8662-4f8f-9dd9-28b8f22266b8.png","iconPic":"5107842f-df24-4ed4-8dc8-476b8a0f3ddf.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.11024","numDisplayRows":"7.87402","pins":[{"uniquePinIdString":"0","positionMil":"752.23425,54.15041","isAnchorPin":true,"label":"+VCC"},{"uniquePinIdString":"1","positionMil":"851.78031,51.38547","isAnchorPin":false,"label":"Trigger"},{"uniquePinIdString":"2","positionMil":"951.32638,56.91575","isAnchorPin":false,"label":"Echo"},{"uniquePinIdString":"3","positionMil":"1059.16772,51.38543","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"I2C LCD 16x2 Screen","category":["User Defined"],"id":"12011600-a4b1-4790-940a-709c15856539","userDefined":true,"subtypeDescription":"","subtypePic":"04d2d11f-9dbd-4a2c-b6c9-835d97151b37.png","pinInfo":{"numDisplayCols":"31.49606","numDisplayRows":"14.17323","pins":[{"uniquePinIdString":"0","positionMil":"-26.82198,903.07729","isAnchorPin":true,"label":"SCL"},{"uniquePinIdString":"1","positionMil":"-26.82198,1003.07729","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"2","positionMil":"-26.82198,1103.07729","isAnchorPin":false,"label":"VCC (5V)"},{"uniquePinIdString":"3","positionMil":"-26.82198,1203.07729","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"273.17802,1353.07729","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"5","positionMil":"373.17802,1353.07729","isAnchorPin":false,"label":"VDD"},{"uniquePinIdString":"6","positionMil":"473.17802,1353.07729","isAnchorPin":false,"label":"VO"},{"uniquePinIdString":"7","positionMil":"573.17802,1353.07729","isAnchorPin":false,"label":"RS"},{"uniquePinIdString":"8","positionMil":"673.17802,1353.07729","isAnchorPin":false,"label":"RW"},{"uniquePinIdString":"9","positionMil":"773.17802,1353.07729","isAnchorPin":false,"label":"E"},{"uniquePinIdString":"10","positionMil":"873.17802,1353.07729","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"11","positionMil":"973.17802,1353.07729","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"12","positionMil":"1073.17802,1353.07729","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"13","positionMil":"1173.17802,1353.07729","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"14","positionMil":"1273.17802,1353.07729","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"15","positionMil":"1373.17802,1353.07729","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"16","positionMil":"1473.17802,1353.07729","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"17","positionMil":"1573.17802,1353.07729","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"18","positionMil":"1673.17802,1353.07729","isAnchorPin":false,"label":"BLA"},{"uniquePinIdString":"19","positionMil":"1773.17802,1353.07729","isAnchorPin":false,"label":"BLK"}],"pinType":"wired"},"properties":[],"iconPic":"d8a1d1b0-d05e-462a-97fe-7e9bb74087a2.png","componentVersion":1,"imageLocation":"local_cache"}]}PK
     ąnY               images/PK
     ąnY�m�ځ ځ /   images/1c49e1bc-8662-4f8f-9dd9-28b8f22266b8.png�PNG

   IHDR  �      3R�  iCCPICC Profile  x�c``\���[�$����WR����~���A���A��21���1 ��'�v�.��b p��'�@�\PTt�.��;�):
����!�;	V�d� ��H�$$6�.`M6J�DvHriQ�)ħO2'�N����&`/(m��Qs����$7���ط�U��gլ��_{��K���KR+J@���@a�6��E_�' Ēf20loe`���SY��������< ��Mۋ�l�   	pHYs     ��  ��IDATx��Y�egv��p���s���f��Vw{��r	�[�P�H^(��짼�E��y!�8	� Jˉe[R"7�I-�MwK$�IY�t�{�aַ�����[��$���s�>{���������O��?=�t�׺������g����5|��t^���+�����1�����k;��J��_��7��I�=::�����>�x�{;����_�qx����<�+'�	�}B�������~+��>�K���4y�l�o��Q���'���@�A�kk?���Wz+����]J	���GW�Ի�P�������k���V��ϟ�͎��ѷ�h;+���}�1=���j�����Or����=/���(�^M�<�#?�Io��M��������o���� ������������<a*'1��&r�����|>��lF�f��Z�L�ɹ�t���k�n�;��n��gN��a�9�ϵY����c��o�'���7�����T���[���1frx0�fRs���z��7:�ƍ�p�e?�nԚ�|��m�I�
3W�j��ͼ}�sEW���}��xc��=����4Id�y^_ot^s��/s{�ر�M��Z��/EQL<ϔ���n�����_�w��W����key|��\����ҏ�}G�M��y��-��}��}�T�w_�Uo�'s��v��=�πi�({�>R�*=V�
?0e�Z�U�U�ǀG;�6�%N�Wz���l�|nG�������O9�<��M�?���[��S���'�"��8�q#�#G��������!��[�M��������<f=����5o�?�6~C�[�V��e4���n���k�s\������d*�[�V��y<J�D��$��3ӽ�}���(�zog��~�=>�~�s��~���h1����?|}�W��h4�=����♳������2Wn�@;Ӄ���ζ�!h��T�5��r}�N��(0UҌ�K�	Hu�;��!��? /+� �/�2"6)���{f�$9����X
��0��G:n�m��I��h��G���e�I��K��x��=����@y�vV?=cy��^�f�Za���y��oL�8��]<�cy��h&��z�q���/�V��kv���H֜����7o�:�ׁ�1_Ij�^�yJ��;�@9�M��]����Sj����^g˳}+,K��DyZ�k��q��x!߼���-�z��b:x	<F�Lo����n��`�@2
@SB;��@s&���������~=(L�k�I_&e"��W��.��8dA�6���x@��&w�5�ȍ���km�Ӕ�PrS�#M�k��Ud���&fbM-�&�D��@�X��๡�łA�D��;�[�ٕ�G�/�N�wS�DE ���wD��̄�n�^����qk��x�1�B�03�|L������4�q�;����Ad�!�����ڈ,^&P����R�E��"�H=a����Y��b]�*�k�Vc��z#��н�B���U������g|;�]�YH�,�٪S��Xֹ T�}���}��H)!��9���v,�c@�{�֨S�F4��H��nvVi�v�
8M�C��Z�����Ծ�i��q�pb�J-c��|f�^p5��o��ͷ ֘�^^,җ��"e�<!��ID��ޣۇ���u� ���H��L^�Y�e���wdN�w���N���h8���A� �Z�����v��?�! K�QW�i��Ç
N��/}�����D���A��$�xy�#3H�KH�	l1_��?�:�.\⹙����x�f��F��9�\�/D����׵V
!a�h5�A����T	}�����~y3�ZX�s����h����3��L�7��XT��/�(R����������K�|U����0|���w��Jw�ģ��MFW��Z�_��A#vخ�w�g��\��^�Wo��^�a���I�TՇ;33Nk�h2�ǏF� TIJ��XKGL|x4շ elO�<>2��Y`�O/�Ǔ�|y�q���j4J����a���S'��˱G�#S�՞�V��(ؘ�4�k�m�ߏ�A�b�`e)�9~�[�ȟ��5��oc�x�}�W�s�w^�/3+{���5<w�0/�7SUP�c.�<Zx]��U/"c�ǃ׿{O�6�^�{����@�vs*�+0��k^����v�'L2��@�Sx����Ǚ<U�}_���'��U�_���C<�T���s���+Rתo��2m����ߕOY���U�d
�R�K�|�Ș�Y)��	��`-@�X�����eO�o��)R+�<Q���B�;��[~��/-uWW�7��O{�Nq$�P�qtthے�{�cV�|Y���:������S����~�ν��ĩO+�|�A��Xh�Uyy�K�}�j��|��:��g8�z�)8<�gA�, l�H�=kr2� ؘ����Cs�lqo������q�ټʌ�U������j�&5�5�1A��j�S�����M��}��r.��)�}���_��x��:�7F��I�,0��@&���I�t�q�xr����S��$���ϓ��0�'�s���X$U�S��Ju��9?f{6�1D�� �v��`�'��Uf�W�i����% �����W02�4f�M�X�Lx���v0��p6���7�	/�*�����4Mh2����o(H͘��R��b�8L�3�[h��(��h;��a_�����E�ǈ9=�J��1�:��*��K�/38����nF#"n�grlm����`m+�l�s2� S�� �*�2�ʂ+e�� �Ff��]D���
�9�[�&A�:V��m��]D����?}���v�-�X<0�T`F��C��?�g������W�a���/ ���I4�����`���X-n�Z&(Qz����s�Ւ�;	#І���3����)k�ܗ�Q|k���t<���l"�����	_������1�uVZ�vA[�5V�ĺ�j��:?���N�06L�/9� mԱN�.��;�1��nu�ϢS��S���F� mmm�?'���$@�Z�ۢ����2�e�Ӑy��##\�5$J$ϣ��1�$g��wg%Z�K�r�k�mU�/�d���q+��O�����|m�ߵ��� ��x,4-f�����^m��ќi&NB�����z������7��?��$Y���O�:�i�!��b��@�euu��J��޽K��{���"�<WP������Cz�� {U*G�z4�}���W���R� 8J��l�[2.��9u�-��K(� ��zE�"ڢk4�ʂ�;����������ߓ���~�����:OvYC�w�NAI/Z�![���ｏ����뇔s	��Y����H�N�����;2,#^���k��}V�������,��_����=���?����;ߓ�����?���h�+�k��X��Ԃ�x�hʴ���4����4*��,��R{�8*}�����f�&�J'�}x'��������,+��0�����ͅX����Xx����P�T����d`+�֥*����D>��e~��@=R���oC2�݈�q�P�p��{��n�,��~\A�d^��Z���
���3������|���@ͼ��B�����	+�sy>�Ё���M^g^�c:w���wx�v��SMXִ�瞣;���p�����jf�H��0[�sYރ6R�-�^^�౭GS���%�_|��y3�Wp�|���t��.�#&��u���9θ�@��$ ��� ��@�I�E�N�LX����u8�(&B�|�L�@j��BM��`�"�(�x��Dk���Ӷ��'j�wn)S�$���v3cQ� 3z�@��.��2�J�3jVCr@�Ʒ�
�*���m1�l՛ԬԄ��m?�\A��Qy��})ϓ�B�s��G��<����v��x�`bE� �X�I\A���{>ڜ��f ��#�ЪZ-��bl����5�����b����	y���	��}H?z�/�����0^��u#v������`�QA�gs�K�T�Å�x��:�X�ΊK�X��Eg�8�JsF�B(v|�D�nJsW�0,L��z���j�i�k�������q�<6s�%�����I��ꉻ�1+��였�T�{��^��<�5Vc�3ap͚���3�]�g�aU�Y�I$Z=\�+�h�P ���t�x ���ui|�2�a��S-b�c!oXz����F3QP��Lf��m֬������G�ӕ�c��-k|��.i�a�>�@�l>��3��b:!`{��)�<��P\w��h,�.5�EЇ�n^�k�⫠sʟ�O�|}�r� :����r���@XCp �����d4`Ņ����@���w�h>b�Ia�,�/�@�e�����4�-�����*���2�v�c| 2D�Oɼ�XUt�$������N���QLԓ��;�2� ����ʛ�s$�����T�W;�S�A-V*¿����p�k2�?Phך��P<�>QQ5�V딇5��y�T!����� �Q�ώ�`��5�A���,_��jP�|�����e-UE�2r�3n�X(]�v~��ku���<�,�����#�;�>�U��a��t�
0� t
^���ђe� ������I�C��jn�����)P�;�wX�6b��0�-���g�UB��*w-���+�#
� ҹ�Ŝ�DAY�W,m�3�F������,�F ��4��3$cdd|��%1[��z�B	Iԛ�&��-���z;�>q=x�W���~D�̈�5�<#�+�����`_��iq��4>0��R��.�ݧ	���8���G���R��/U��rT���04p�#?�!�8�q�Np�����>k�־�n�<��(�6	6��4���*a�R�h���+7���f�����`� �&eXAU>�� ��,��0�v��G�R�"�ח~�j^�2��b��7���D�±a�Q�	`	��w{��;�E<�-x��ֺ/�.�D�L`qq��h�_��]^��R�X$��ќ	Ze2�k��5�ˀ���a�A�*�X��ł$h�sS��9,y�&�
������)�ׄ��7IY�mU/`�TBC���� #���L..8����-��l������3��0?�zC-�$�}Z���,��H��	�r���x9X�������hl/Ԗ�Tׁ��UЊ�[? <˴�G�`b��]F��'��EF]m �BG��t��8�Z��@�[��@&�ȘH�Oj}!�<MU9A+.^��S�x�#�H�w�Kx ��h��(�Q�xK������4��:�F��stvk�����i3Sfd��)(���4W͜I����x(����z��vD��z��
B������"`��+$_�Z��j�	��kX���3�D��r�b�X�+�!B8���v-����Ġ)�[Y�v��d�۬�ba�v{���T̠�f��XglȊ��HXK���	�)���Jb�Y�f�-_�"xq`\bjy��?G���g�S繬�v�yj�����7���]:��F�_~H�ޣ�z4�ӄǽ��k�u	ߘ�܍fP����AM�m{����>?!x��|��P�3��y����3-Q� 2p<&#�pp#�6�V#�Z|��̦аx�����ZkjRk,2e
�&l�� �P��3e�g|V��vܵ]��I)�0xNB���oFA���!��FkV��G�Sa��R\W�9g�<͉|�X��E�j�J�������f@���<׷�qX)���^b,	���@>�����3�+�Ջ���R���Z�ߦ�O�����0���ҁ�d�I`�pG��z���!�^�~��7���U���Oԣ�M�@]��M$vЀ�P�`�)BLB�-�.��xxA���n|���9���<�a�f^
�&��؆O�֚���%�FX�-�P޻4��R��x>��̝��)��McK(0�Ҍ�1d9�w8����$<�g����f����&��į�I�xJ_�c�H��	��������h��vA<�v��є�����]:�f���]������F��0�4�S�g�`"c��1�vAb a� @�B���B*�[`i��X8_�)k��!\惩,80Nc-+`�ά��*��p�Ohk�jl��K��B2<`+&Р_U1�K�����,V�=�+��9�u��_]���#�����0�FG,-Hn�q��0���j9	��ꉬiB�$�(c,2��W׭�&�puɕI,�����{�`^�d+Ѐ�D�x>�͆,jX�b!-O��F֒��X��T�%�(׺ETxb� G; �"���V�Ո�*� �\�����5g���` �Fo�1+���&��
(D.m7�'��c
��ў>w�����3e�"$��?�h_%^g�
���m�fp�\�|&T0c��$d  �8�
8�c�B;�<(K��k��!��D<��� }^S���9�c�#ԫ��'�f�J�)���/N�����z��y�hth��e�m[Li>:Kr̔�������y�a��P�2�}����O��6�� ��X7X�����ź3(쮴s˸u�8��Z"�/M�֥7YZ˚عCH���R�s%P,:�`MF�XE�����񋅓��yX��>X{S-KG��m�}�{��Z7$,��*l��H_`E�d�&G�hܪ�Z,�Ti��PYߞQ���h3����ǀ� �����)z���t�	�,�n=أ7���{�.m�i��08���XG�]�(1 ,=�i��?mNY	���=���<VU몔1��l�� �!�H�3����X��F?�:���p0�����X�b���X�[}h�%��_<�?YX��[�^��`�&��@���S҄�@�A����]�sqT�a�,�������Xd���,'�:j�`^�|��^�<+�q(�i�uV�!�	�)�k����2s����;�Ij�> 4��,�5�R(/�⹉�=���t�Ԫ*��(Δ��?O�n��
��N��%ԃi��b��h�5Y�1<p��#�u�$�t,��@@�E�ސ��p&C�x&�U�w��F��#�'��2 �B����4�0,�aY����B��%3��X������p����0��y���w*y ��T1dE��aʓ�R_�F����s�w��ޮ��[{��_�'�o���K��	�0n O!�I�����0#D�����������Z#O�1�˱�$�O<�k�"I�'�`��0�u��83˂��rc#p�ւ6�D&���Aᜅӈ`���]��W��/���b�k`Ń��FMXx$�-�,6@՞@����Gk� ��K�*�e`->+ř@��D�X��u�|! �9�u:p2e&�-��c� gε���.���W�D��F���g-Lb��t�D�SNLy܌��5��L�x"!΂;}Y,��<u+������a��,t|�	LB�3ށ�D&�|ƛ*��m���^��R�%!�i,��d������ ]�T"�����ɥ ��^L��1;��
	A0�6����$Fp�U���f��9熅�x8� �`��!/���A�Q�@@�{<W���,�8�?�I�@�$~V2x��jT)��
�?J$�(���N�M�w}a����Ӆ�@b�Y�
�,�� ��?<�O!4���#j�s�O�i��.���'��箜�+�N3(���M��4`:�e��
�6	��"�L2ik���q�y��d��e��uVF+���) �5���X�JC�҈/�0��VK,ryv�&�@��u2��ʪ0�4u�@2�7�ܡh��V�8�Z+����[������E4K.�кky"��N���WT�Zh�9@s���7�E�I	5���e5�!q�;�`�k�_�x�z+��G]�ǐ4N����=��!���I[�l��?O�/Л�O���tgg��
���*�<��H�"�i�ڦ��DRa � e�V8��j�%<3݂'qQ�I�A���Ա���f����"�ǭ�G����b�n�%����J�M�@PA�c��>J�a��\j^��%�+d��#2��1y������9����Z�|����L=�ܤ�C�O!��^]af}$q�]Ȇ��b��d6����R�
���`C�5�e^P����Td�z4� Q���5�Z�B��"t����q�`�7>�6�#rC���!y�eF%���^�zF��h��i�ʔ�9P��^�!��2��7C�n �ڬg�+g��@�?Ǚ�<]]��j���u�Gƹ�+������P	
�[ބ.�_�&�Z����EA�ϊU�	�SQ�юj��JxϘeN�+��g���
5���v@����zgE��h�՘�����		r�.2,D�ð�5�ã;6G��v�M�	�!�|Ɗ��,��V�����ea" =�`G��k�(���LL)�y�ZQ��d&�+T��y ���ɨ��U\�4�.$(JyBa󬬰�`��H��0�h���A��cAX���L�05�Ժ���.��2`A��)\�M��H�?�z���h���̝�C�����	[�K�1OW� ���R�`2B���qr���� ��X�|�5R��,&^�6*(��s��~Ɛ�DCug\�_��
�g~��τh��8�^��_�J�?��[h�-��}ux);27�jZ�f=/�`4���>'�Օ��U�,J�ϱ�Bg�=uɇIl�����eؑƟe��=`���,Ɓ��ǳt�5<LKnhGz��ui���T3� �^��I�T���_�
��63ZV,ތ�����s/<G癱�Ɉ���|2�n���P�L��E"�H$X[_���^�-�֪$(Ur7��3D�Hr����%#X�,�;�1����Hc����X3jk�$-���0��`Occ%y�ę�[�5�||!T��5�0�g�Y�
Q�$�\3��i�a^���'�HFg�k0�5����Zqaiu�u��p�/�H��ә��@�G�]�����w��r�Xِ}K�V� ��\7�gs�.ܿ���=Z�S�ަϞ^�n�9z��譻hJ�X{�����Uy|Y �$���?�ޟ�ņ�T�(��[+�K&p�%���a9YF!��m���d#|�S����VKg���W���˂Z�@t�_�:ws�Zn���x_Z�� 3�{�oc�H[Z�2������E^��e�4�x�`V�>�YY���$c7X*&7<H�LU+����x��,W��hH��}���/�qrc�ɮT�\�j��.�i�7xU�g�|r�e�A\V��*���x�-�k=�H&~Z���g>n�%� [�s�F��$4����ǁ�B���Β����5�����Mx�|6�dG�2�̰OW.^�3�+���M�rn�1���W��gr�S�&)}p�޺~����F-^} O�1[苡'b巁8s�P~�C1O���P�(H�E&Mļ� �|��ۦ�$h|�[	Lڴ�FX�5F��������tjk�r*��0�B���`D�"�n=:�ݣC�Z�N{��+�H_Ժ���ŀ <�u��VK��^�djAGj���������d'H��q�����Z���|e`NkE)A�}&��Q�iJ@�+I�� `�2PL��ȁE�N���G��u� �t�'��e�m�i�h5��N���t`*A�{bǑ����o�4]��l�b��j��9S�4�r^!�Ǚ�m��	XZ�m�z�g� ���R��"x��La�9�}{��������%�Y�=����|�G���0~l�Zߩ.g��*b?��D�]tey%�������Ba�ecR���\�iLk��R���^�������P8���}
X郓��n��y�+�kc����=���6�HK����?�M㙍IT�l2A�C��$�nŢ�WJ�C_CAZ��4��B!��=[S�
�2����`)D�Κ�q����D�G�t�.ֺ�qؐ��Z@_�X��Biu1�\�;ۏh:��0x1D	9�X<-���:���l��[:��pk�����j^�)�FM��cn%��<�r	�[ G^���i:��р��$�nOڵ}��Y�w����/޿C��-y�j��v1��P,���"���)G��o+��
��2�l((_'f���ʍd�X�
��BԮ;�e��W�j\<*�}Gq=-{Z��~��<X��=���Ci�uaf�2�~I^�'��5b}�f������yvE�N�[D�8�X䃃�<SK������L�h�zb�S?&u�yV�fZ�r�����v�����k���oxvl��؟3a�SSnپ(#��zfJe�L>֑��:��a=����c�BBb*Uʉ��~+������[�K�%֛�r;�>;�gk�Y�T��1ٓ��qm](
����:5$�0���7����3OQ
�|@5^��t�<r.I88P«Ì�֩��sW�������G�揯����Y��gp�k%���"1M�"���.�?��ƖIR�e<P֢�:f�v��vUʑ�t� �2#[�t����.P�ۢ!�]ڗ8т��7�U��B�̅s��?�����`��5��/.��w������Y�g�:&Y-'b��z�b_�bѼ���+�-�5�sM�@V;��vb��?+~��5k�Il	efxc����%Dc�ڈWp98���ض�&/6;R2K��ϑF�v[��ک5�lZpֲ����A���c�/�4kc�~�\Zߗ���6�3�]-R�4S��;~�l�Ɨ�j��AkD"����9	���"�,��$I�<�b�$�.����`]��
�by�T�Z����c��X^�Qo�ᦉW�4V*!W�o9�ڳڭ_�;\Ҍ�J�Yl����p�k$������Pt�C��p�~���yZa���{�YkE�fT���ڬ`5Y���e�u��-(������)@�)��ܖ���u��L,"�gE�MU�op��b!� Z`�I���({�8RX�`9��H�0��L�Yظ@h8i�I�bKf� �zVA��O�|X]����Ʊ���8׳-��hJ��\�{�J�$�$�>�Lw	ķ	H�E���`��%:�5�U`�e�#ㅶHVjg�YUJ`�j!�Q�zk+җ��-:������٥}V����x@g�+�{�ɪ��������
���B�"���?x\�)��=
V�d���������Z{�H�>�2 ��n�.�Xc��G�2�2�Z�<+�L�u���)�䶲��,�(�(�,� D-3����$^��`̀<�1�(��p w�1�׵T� �_3�mj�J���$��H�-��B+>4~��$Fc���"���]��M����e�lbr�_,����{I����()����br�.r�Klf��c��k�F�!X�ۙU7��Ce��W���0*���/�ā8���%^^h�@��%�1�ĲK�i���uMr�)�ruVM4e���/��gϯӗ_x�֛��#J����U^�nK=�B�HEXrj��֘�����t��i�ο�3�?��ʊ3,��w���X8c�Y��\[]�x6�ߛoz ���hAH��6:��#�$�I���Zy��}���U����<A_�t�VX"S�[�i�ײ1(�Y28D�}��&\ ��0������{��O~�#�����0�oр���A�$�V\:ab�ᨹ����R���#[ r�i���vW�2&(���q("���%ط*�U�JV��p�,Y�a���M�	u>L�T��M�"�� #cr�A�Z��J����ܝ�1r��hAQ�pax��N���}r��扫i<���sY��j���ϖ_�E9����?s)�*�Qb�0E��l�:.a�}
�MM�l߄���Z��]�/L·u��{�N�3�LI�πXRhu���B����z�eɺ�琸��4O^B���|�0�o���.�H�5!�@��K>fcM 9��-=儣瀬������HV��MM�S����Mj�1���/�W�����86Z���)���xFrZ]����J�!�yH��>3�C���f��v���K@ mo��f��
���r68fc��3z�A}B���~�%�|��Pceu��?;�~+�j���9�[���CBPq�ۀk]��o%L� lʡ���hP�{̒�븵���3ZZE�-��Q_�ǀ"^4a^���	���R�se�G�y[��}��j�w���;4B�8�9 �m��xq�ήu�{o��~p�>�W7i�-�J��#)we��퐨�2�_��R�ķ��W���[�B���oiVʨ8�š9ԖCM�l>˱�T���s�L���_�>�g� �{m�NR�٪J��g���Y{�S����
�J,�EK���U:($�9:GW���t����%��W�5:��&��JNPtA���Y�&CnH(��EBU��؂$;7~�n�\�1B�%APB���W�`X0
�}Q��2�����W�f��|A+h���OvN�@O�����Xͬ���}�	s�"-Zh}�S�����c�{$l�W7{$'"q��h��{P+���|�)�����F���`O�����Ym��mR����H�X�U�4%޸b�e������x���������R��VC+=z�'�Uees�W��0d����h�!4l]�Ccj��c���`@sf�n�*��/}�*}��Y�m?������M��x�����d]��ۍ�kp5M&c��|��C����Vi�}�?�Mo�ݦ��H��%�J�(� #�L�Y��%,��,�$­6�yDC���;�<Xa�K��稳u���`D��[ ������R$`����[(Q8&b�~.#Z��P�5!�-W0�1����� �R	"k����\��]˵�d������e�Cژh�I�8�Y ��D`����x�L[�t��=�B.��e�c�J��2�0�yR�Q&�ei�lAg�+,7?����PY�}���vjA���gu���ˆV�A����#�����?�EǏ"�f�sEK��kA�곥�mʊ�GuI�Re6�_}��k��B����ʝ��A�u{]Z�mH����mn����ɷk�x� ��c��%\j�%��֊(g��O�k?NlU,�j�F(xU$G�^&�ʖ����;�;N�rnL��\�[K�(��ɥ�spmZ����' Z��h�K�@1ɵż�D6������k���ɍv����u����?�~M�Z� ���6�oAco,���lK�Q��BMXy~o�:`����X��gLh��y��t4�̓Cj4WYih�bO��K�l]g�H����4~y'���c��Y�.Y���_�t��S�xo�[�q�-Ą{�\^Q�}+(�K��xR��ue-�>���`�1XR�ą!	���ƸxQ�}�t.����<&�d1�[=�c��Ͼ)*ٸd��x�<i��;�h�4��2P/ޗ�%z+H�����C�Ǐ�l>J��{�x)������ۙΩ� ��/~�~�K�R���t�O�*5YѮ��ެ��/֩���x�6O୙ͮ!��c��"JFJY�m���A�t?�Oy��b���4��xD�����Vo\��iJ�oczb��4dm�[1��H��E�/~��^�@�L�c����-�n~��j�&�f�uQ����xwuœ؝j�ܹwW�VX��V��wĥK0|���(���5wW���{dAb��ֲR���#3S�'��jb�d�֩��J-�v ��=���}N�9jb�u�Pf
�=!�� �^������b�#GK��
D��a��3�4'�X�m��P� �Qtser���3i V:IZ��>c�C|�]ஹPLJm�mbP��i�VJY�F���(Rn	s=��R-~�Ql~����$�p[�AP�	%+&YX��V@/���2�t�BX�
y�ԇ>jq�M���JX�r�".O �)�����ZG)^�9�I��"p�L���b��TF(�Q��)�NFC�zj`]F3�}p�~�[��m{4���mܧ��T*l�������=	Ѹ���g?�4E|�b2�[��g�����8�P�kC^���B��Z��B,il5rX���Y��}��ci��Z+5K>pb�"���E�#�ܥ��B��q\J����� ���r�)K�[��`�����gV�b_���!�<]���j����$����:�8+u�>��yB�oߦ���tc)���RZ��>O�~�`q$��8�7��~*%��`ρcѕ��@�IIk�Q�$�]���>:nQ,*���S,�~�gz�Ўcoʓݲ�����0餧x���>c�2H�m��кX�l��ʋX�L3��CG�vD�Z�3ZOc� �����Ӻ�j��G	�|��>�ye4����gJd���J��@�"��O���d�i�͵���8�^>�w;���ғ�ݍ}���K� �	K���8Z����c���f��zpk��x>����[��׿�UZ�D�Ἱy
��j��b�o��<ih��
<�&��^�Y��k�h�%n�z�}��������&�S�Xb�_�v��=�rj�X��F���P�,���f�:QQ�N�B�ʳW��'/P�����ԅovV�/����lL�`{?������={��t:W���?|��Og����Oќ��ۇv��q���2�YV�X�.X�_Y��z�D�Ӗm�^YH��H� �X�6�qDv��"W���m+�@�<��8Du��qA��A�����Ai�u�K�4M��Y���X��4$F�� ��=�ª�~�X[�?jB�%��ϣ�}`Q.��ܞ��
�ӁX�4��(��P>��krׁ[��u @n��\-�Z���F� E���+�+�3���0�K�o�n���^���v�(��8�Q��j]Ly��ܚ�f��;�sD��^͕��kǳHWV�Y��\�;�.���74��T�U(��n������������L�׺�����0uk+=z���ӈ���?�S�y�s?�t�+�?:���(��ܰ;#�c�x�����6W����Ĕr6�g��8+J���GĐs-f��C�,@
IPE�c\�Z?Q�>x���|�b�x9�,�*��C�|߹¬�����l��:��]��&���w����pG)/_]��g�k-����oݹC��{��`���>GϞ�>���޻M�vE�k���/|����E;�RL�H�Pj�a��3����.B���H�>���������q��d�y,�w,��O&ֶԔ,�Y5�eK�	�v�k�-}����6v-�N��ѣ��XF]�W7�]���oA_�~NWr G<����+��6�+9�,u���;OR�%9��Vٳ�>�_t3	�Ԫ���0�W�,��XJ/�zUM^�?�*�c�	<5�p��O:�
&��c�dr�_���JyL��<�R�
z��Y�4��[���5)c��t�<��S+�]P��eb�0��z]YI������ٵޣ�j�^|�iz�'��ۈ�-��<Cw�=��sO�P^�e;�^����\�6K�Ϟ٤o|�
����J�g6�U���[���b:|gN���ʜ�����n�m���������מ}������p΃� rOJ1�n, [{!3Qk6�C-�D��th��+ōeK�z�:�7l���Ę �G�j��%�q ���-��R6�2I���-b��A�f����L�8 �j�}�iu��儂��l�;3��T��ع��
���
���~'��͑l��p	0Gm�d.��
��*F偘(��L��"T���.q)VD���|K$�;�8+���c�h-�P��¢���[�AT�`;��fg�����E^�)MY�.8��H=Ƹ5.{p��[f�.Iɲ�ϓ��v4��� v�B!R� 酩�z#�
��W� yumEv��N]�ϖ��퍙;�"�,�4gB�����!N�4G� ��O��X��:����ϡ/5��!��!��>����[�̩޻A5�$��:sj��~�y�_����I���wU�n^W�r���h���2�qH-�T�!alaw,@�
Fg кVs�m߹f��,Yz��h{E��>�b�8ͽ�;ĆJ���uK��*b2��j���Z�Y����l��D"I��<�c�e:N�r_5��y)<�7b	l����V9��f\	E���z2�Ѓ7h��Kg/]�>�m�ڠ7�����g/�}j6��K��%����H���$fE��rg�&}�m��>��XВ�1g��y�UleKP�el���^륣�-�V5��J��L��Jm�\��� ��L^ɗ�δe�퇣[S��e�����c�{$r���*Y����REQ}5��O����\Q����d�4~F�5��	!$�7�*v|�d�� ;�;a^,��Ī�߾�1�1��tC_É�Y�d=��rAEy0�M�uR:�ռ���u�Q~r�gj�q?�|P!���>n?(��/Y�uO��&��?�]k�{V�d���[�$�Ê߅�Xچ���o�7V�g��<5y��+���H���ͩ�4��dE�2��
$3���5n`�H���l�a>�Ʃv����J�ޑ̟	us�F-q�P�"6ӖR����M�e3�xj��9���-�z=+�Γ�V��,&/=A�;>OEː�e"9��Gáy�DϜ=E��=C�|@�پ�%���jsl--�YMI����L�/;��>�;  ��	1:I�%nmX�O��tfu���=��Bք��r�2W&�ɶ<�j����u�&��m C��!���j��Va�%�m�0�oK=ȩ���$l�����Z��&jbΨ�Ψ�Շ-��xw$�@�s���:����^a`Vi���]���la�٤��e�M�eO���M��o)�&�߱5�l�0������@vS@�Il�W�3\���0�(��Ь"��B���x�լ�e�`[М�<��Q9�b\
 ³`鷺�jP��r��F(N�P��K�(S�!)ץ�Vi�Ԗl����ò��(́%�Y%raR,�Qj����n��y�Y��a��~�Iz���
w��Ƌ���:�|�-�|���������h:<`� z�g�g�����?��I�Noү�{G�n޻%�:�*�ݓUѽc���ւ�(�tq����k����O�n��9������d�F?�i̶,��B�6�rZpϗ�o���˶>�w*X餪��2��p4���V�N�F[j1޻}��>Ϟ=M���e��?�c������S����C:}�}�O��=:�I:s�I�0����[��4�g6�p�39���M���Ku��I=JߙGvy�#k�m<Ƙ��`���H���>a�e��';\��2`,Z�<Ʌ)d�*	��a�����Ogi����
h�*�(ڍ:��U^�bP�VC(��|Bf>P4�M��Þ���ض�Y�p��v�(��9X+m�G)p�m�b�P���*���6�%$�m��(a*���؝S�
���D,�rq�9D���<�T��e�)с;�D���95.��Nb=��t�v`����d:����jj���y)�l�R=�2����2�{��M"���Qd�?|@�N���>s�,=<��;P��f7���Ew��+�n�����u���-�r�u[u����q�5G��p{3C����ly4����/�ڤ��G4i-�ZzR���4�,)hP�B��lؠ���[m��j�՛Z���%)U�V1�Z�����-�	��Y���5q�F�_s�L��Lj��x�h�}�lpH1##�H��lŀ=f����n����aGlÄ�p�yDa�@�� ��+��j����^�z�.��t�d�n ��k�����eHֳ�s�ۂ��h7����nt)��E~� �MR��:��{4�b�>�����'��&������B��/F3�:?/b�7�&ט%��Z�+;���g�˒B�>-d��8_�u�5[l�U��x�7ǩ�e�z�0e����GR��r��4R��ufVK�d���昛�"��}���W���
�irg�<�����Wh�Q�7��8�Z�C[�л�������q���w�.�����������B�ڶ%]hɵ��y�G#�·�62I����0o�~�!���<���!�/�.Z"?�!n���łf������-��=���с���r�1��Q��ǵݹ�u�t�Z 
��m6�4Fr�G4����g��/}�k���[��7��ŋt�D�{-V$Ѯ]YG�Μ:M����w)�3���(K/2���ɭ��Un�K��;aV�8��W8k�j�-��I�d����-���ІL�\��[N@<~�`:�F�ؤe��PlC�l��FAjVZ����&]xB��o�@6$��$��@"���*��|0]��a��[�Օ�3[�� D�v�;��!��84�d�	�r�.�Z��N��MfM-�avP�L�0(�$F�e �IϞ���}��;e�+����������`y�n��B��·�DKe�u�}.y��q��uO6��w��T��
��Gj�
u�D��r���V���&���b~)t
G ��,��h�LO�AA�B͕�a��ڃʋ�t���+`׫��ۨ�c��쪀m���lFA���V��=�̀��gok���a��SJO��
D*��&b�q�jͰ����ƴ�D{vc��ǻ4��TR/�5Fy��s�o4�+��Bقiuu��|r�B���U�@�2c�Yt��U��`'�(g:N+(��3yj�R�A!�d���9���M}����wc���
7���2%-H98ܕ"��А
�1�3���ޚ|���k��jѕsg���S���G��@q�U���	I]���A��{R�,�,a�a��RVc��d�bP���T����ֻ�6�;&X<���V�,�F Gf$�)=�;��ww�����`rJ����\Tg-������B�,$G, Xж>�Ժ�VnA%�i�N� G�ѩ�Y�7 ��Fvi��TO->*Z���=I~-�=�K��jq'���H�c�ޏ����7/F�~�L��ǲ�Hi�jm1�gfq��:�;�ڬ0���s�%�˿��io{��{�-�����ٓ��
�:+)�����p��-U8�J�P�w�Ң��۱2�D'�,n[���g�4�q��hMUk���e��e��a�@�*������ٗD�o��k���~��l���5%�[z��t���sO?O#�4�ü����:�<�KT����R!6o)v���S'O���BjU9>9��uc�	������5�@J�M��<���b%�}wZ�j�ֽƟ{9
�Q�p�X�=y~R�!�`V(Z��w�ٗ}��S�&M�l�`Y	Kbou�6�֥T�/;�h�Qs�m�|�*���HS*�w��X9-�~4��6{����>͙6��g�x�+��C Fw���P�>�d�2�� F"��` �D"��Y�o�bxjPHI�9u�,�x�	��>q�=ކ�~YV~]�W9�>��A��@��DE��+�7��J�5��E؞XLKQ�2�X��dH\�aQ�m+�I�Y_;uv����?�.Ɯ͍=�Ed�%ja������D�R�h�Fn�*��sݦh!�N��U	^giD�V��32wE��^|g�Z��4�rQ�^����)���П߽I}h��ԯqY�d����?���9` I�8�,�;��m�x�??��nH��w2�*H˱��)�|&�Z��yDY�,��Z�~ �W��.B�،��to�|^�]�H�b���v�DP")?�@>a��A��+�[[�sgNѓ/K���n�6W�D��F�:>XPs�򆃉���6PlU�-s�)�{����n�C�5J�m���8���@Y<��g0��E�qz[���~�ع.l�ծ�Zg��؜��9�;�KJ�slJo������!������h؏�z<�	�q	�0�1Gآ,Fm̖�O�˅-l,VkO3�*���gWU�)[Ho� x�Pa�J��-h�
.HyF��3��n4Z�Ecn���k�E�2����>4sxI�-��i~�D�y,IH]�A`DV�F����Y����3��y����x�b��;?`P�C���Wi�[���6��*�I��Pk(��3��l柋�+��T �w=�r�����J���}��	Ib��/���ŤL��s��N��\T|��XlqGDǘ�Y�t=+���ْ5Z~	X{g�Q�l�)_�d�m0S��Zǘ�ſ��&+ C�զx3��m�}�ߠ���ߦ��]:e��i�/�oݤ���9�) �~�P��ȕB����Cv*Ođ�er���W�q`a4JZ{7�%{Af�̲��O>��/��e��]l��$QxT6�5�ָ����a=�U �ɐv����(m�.9O��SSu�}�=�u�=��"��O��>����K�/Щ�$C0��a=Q�jE�	����Cs������k��Jr�H�+�v׎�;�Ġ0^��Jh��JEeª"C_��!�8S�)5w��MA&����C��l9�7����}���]��P��M���
���(["��,�u�u-���E3�}��9�%�d�y�#�Ʊ'uq�W�2�g��^��HV���%�nK(�⪇�k!���e� D�1�Q���)�� ;Zy��Mݬy�?�R�W�����S�.DΓp��f��k�N��Xj@{�����݇��6f��i>��+��w�=*<�Ϯ<��Cه� �$X�n/nm�&k%�@�W{k hV�������,g'�S'.X	���t��,ҫ띦����yHR�U�-��.1Pm��֍�.��X ��o�<MP�L�%Ss��+;��MJ�:\E��Ơ�ؐ��xOXr�X���.���|e�/X�FS��[uIF�f�"��kw۲��S��ӗ��y:͋��n�Kس�T@��Z�0aTU+C��HV@,��U��Ќ�����}�t�øAP�� \��(�h<���8)+�f#�
L��3�!Xm���/k��l0�I�����zJ�T������S��h>�;��!ݹ�M���m�<�'SI��n=l7�8q�����BK��#��C��Tr!\.�\�jʓKN�YW�}�rs��K6�Y����(�@�P��"����h�.,Rl4���}����H��*�ި��]�|�>��z�Go�lx���\K�u�^�H�@�&N�fz�1Ǯ��>'��U'e&/�b'M�ּLI1�!����=���eO4K@(���qĢa��Q���j��%kg�I�ˏ��/h����ln���;�{�]����K�N�谒�)�������Q`��K1X��h�o� �t�Y��x��Y�� N.��ly�kP�B��Q�]k��i1���A\��[�+�ׄ��p:�t6fPg�ܤ瞠�+t~k���pZj
C�׫Z���%mB�1����aK|�&\�-����H�cO��;�  g9�[�;���[�>E�>3�{��-x/�_Ǭ��z�-qUO������������zpxDs���i"��Yf�3�$=V�ǉ��B���h9��Y�U��5�d�Gǖ�Oi\���ri$�wZ�Y���s.�dD���������� ˅���=na.�v~:w�4}�}D[�uZ�X����Di�m�$+��j�o��5��l�.;_��Ud�,cc�`IJiٕF�G��(
�e�hd?KX�:/6g�Ym-�� ���ط���KF�i��EKu/I��4ll&��AP�V��4s�Qx��_6h��Y��@t�GvB��\�6�1go�����F#Z����?,Y��f]]B͚O�k��ԥ�� �%F�M�m^��Ut;1hj�zM���8b�֏�Qt|�؃P\��I�qY˺U��sI���H2�e�}M� �Z�� b�`763��J��Rk4$�92����xW��AyO�� ��2��5KUb�fQ�	�b7@�L�_�|Y��wszČ��K�oݢ���?ꋵq�ޢ߃�����L$���1��m�U�3dsk�%��\B9!d%-���Os,�����s���Z|F����b)���ER075ط�獁� ������֩-�����������������M�m,�-WQW�����b�	=9	���A��.BN��`��&'��>u����#����8�]6^�YƜ�����ijfy]���V��*�U�T�V|�y�#�x��=궺t��%�{�M�?�	E����x�����w�h�!.,Fm�4[��%0w<�D�g��]���}?�X�0~ܺ\v/+:K���b[���<B�H*փ�I]\�5KX�Z���o�)zU���OBj��6R�jI��q_jcǴ�`�:�PbG/]9CO^�@�y�U�HN�zt�k�g��ֽn1��Bu�������)��4��Z�8FQi>�S�$:��<)�1�_̵�>x��(��������j�A����y�ހ( J�%�]��C�3��9��dF���wtDw�=�{��A���X����[���fb���Ji�py�2�0"���/_RO��\u�r˳���l�w��d�q3:Z
�<G�U�B,��u]����u^W^ �/����M�r�>���M.?��
?�֨� /5d<`ctE���Z|��]�� "[�%Zn�qհ"{�(h&)}��lY���pi7�A�P�Bbk4hn+$��v�b���۱X%�����ʾ��#����O)0N:N��^�dpPK`<�0���Q|x@-�m��x(���[�]�p�>���R������\�!Jޤ��"DB}�$�	"s�#| oRG-����h�"�4�<�:���h�Z��`���>��dF��ga���-j�}j$b�^��.I .��v/��P��8�BO��DEY�}��و�Æ� ���H��X��86t�{��<�A�G�cƐ�[�G�n?���{t{o����[p;��c���B��L|��S[~����6J�J��'7���|��/0��@���ۢl����#N�L� K�I��l1�0����tY�O�cmnnR�i	4��?�s�җ�D5VJ�>3�{�
���G�Z������
(}Lv��[�����,�cY��5?�W��qY��[4�'����Ȏ����2$;��٧������;��������@���[��g��4�5�����/Y������Yem�v>>����ҧ�ە�#x�*,�_�G�C�֚�vk�����@�xM"��\�K�<C_����,˃��!��1#��C~Ɯ��|X=�&�Њ���0�D\�?��_��2�+Z�3��%�(3��3-�]6��=V����p/�D,~�M8�.�/���Lc9T�[�K�_�
՘wW_��B�}���,㦴wpD�ߺC�v���`:�s3��h2��ؒM���)
Ҍ��>�|.�U��"���|�[�GV��c���ܨ�U�N�q�Q^��x1�����s�b�1,&�cJ
7�DC^��wX�W����Ӳ��a4��F�r�l[&0�w:�����r˞��GȥX��un\�g~�^�^E�ncC®{j�N2��V���j����=u�X��:�:A��B
�Eʚ�i�#� א�x"{��]t�]G�F/;5���h�@{��R��x�W��M����L�S��&��Ң��E:s�4]�x��z��fƌ���b�lI�j�e̞���7`���ƃ�d�6�d���"XH;,y9��d� �Ěht������bX%�K�d>� �T�D�;��@e��z��	�Yٰb F6[.�V`<s0=�-�=�:��2�*�3�� ��sUT�\m��艟�J�φt{���{@�\�E?~�� k�;�]]�>��c�4_Dc�;J��,�A��mcѲ d0�η��%~�q�r{�栮Ӕ�|H�����"�BW�F��ڪX��U�+y�Ӧ��4���e�&��#L��-��oܔw?q�2�>���Q�q������D��BT���:r���}J����8!�qq���(���ZB#�(��i��g�V�� �Ǵ_T���{ǀ�G��խ�~ϯ+Z��:.^v	�=v<��R{ă��c��QkI-FT�x����ﬞ9C�g.����ĥ�;|���ᏯS�x�n�i�-Ú�a@�bzKfy����1 ���o�l��$cĒS��\����N�0~T{q��V��Ÿt�ѱh2��Rt|����L _�o�!�m:�"�A��K�7��KO�+�3/R�eI�/n�C���ʈl�xʀ1��`��{M,�T]�v�
���� f�R����.I��yݝm�,�z��`)t
��L����@k�'�>�=M����3�ڝ���o����_�)Z��v%��?�`@����_��й�g)`@x8�҇���{�>�s���x�"�|%Jc�&�*�4��IJj6��p����,�,��_���滸�o�.R�\��quc��L� �R��h a�b�� {FFk�[�?��e�+0x��v���Yo�+�<���(����\U���a�����25w�|��_E������Y��§������	)0���(2R�����<�vk�R+�/���+g��̺T��7so�$Iv��w�="3r�̬}�Zz��Fw���"F4#)=�LO��L2=�L� �ȟ��3EQ�"4��Ah �7��z��=+++��#�]��ν�YK/3/K�Ȍ����=�;�w�?X�P�
mw�?���}u��Jw��D��9rX��xA=�p�!�o���O|� (����wۖ�� �y<���Ӏ- a��m��uǏ5A(1%�����;Ϫ�0��̽³������>S��`50
_�Ť��(���������A����C�F�`������9��a���m9($k�5�Ny���^��0]��<sQ��X�_����z�}Y۾-�|Y�� ]������ a�4���j�d�� :&A��O��������y�4��䞡���R�ǜ� 贤�/Hk���sK�v7��F�̩�0�{�.1��p��\���}グ0�(�:��ƽb6KsϛI��� u�>�:��y�g����x���P�  :�OK���Q��v[�O�șG.P�� Mu]�I���^~C�\����$Fqx�������ꏱy?�*�dǰk��y�t��yy�׭` �)��\7�̔U�#(�ٓi}�Ӌ���Gϝ"FQ�B����B����<`TC��\�5�>�("h�]�~`g(p�"�g0�q���T���;J4Dw|��-:'r��=�i$�|1�@�25��8q)`�nhyͱ��|,���v���c)S�}�́����sI�zUCR����� �T&���n?n�B5'��+��g�a����>�k77e��-ݾ��e�;�jD�[�n���YF��i����!��0���i�C+��8)�B!@E���nC30~���~���A?�|6tʹ�L4=G}W,No�=��+ȹP�����`���p�&-���(3�ì�����aמMW®Z �j�r�oy�F'�&mO1��b��8<Kz6�2����,�Σ8	��W����I��J��(�C^e���|��B�ήt�6eZ���O��o<wQ�{�.�T��7U����W*� �p��kn2��&��6��|������`ݵ�m���ώ����!��\3	�>:t��vg�l]�&0#��P���<�M��/ 9�ט���5�G-�M��d"U�dݹp�q�Ǒ��h=����^�������)l�S��\���T���TG�k{��FE���=$�W��|�[�#�^�_�����$��
j��̊Oc?Q��,
Y$m��وLv,��^ǁm�&=������Mz	��t�����9��r��	+Ա�����!ԗ�����#�[�Ȃ�Ǳ����Oʒ�7�V��#�{�"w|"��)���������CZ,��Z�#�+r��q��@�kR�R����e���m�s}�Q�PB������Ws���9�8��-Kx�=}6=��������6dw��E��@1q�{�� ��,�KN^��H�Q�%
��
rr;]9ztI�T���#'eq�*�S%I����&�r��7����s߁Q�����Ӝ��y�� ��FG�46C�U����U�%�T*���̜��g��:h��X-X������D닣#C�@|
H*:B� ���^�F-s��Ɉu��^L6�u�RR0��Sö^�Ѽ�\C1�fy��F.��J�K��Ҝ�?T�G]���Qи#���ɛ^�w��P٨z��0%�T9i�N�.ښ��':v�+�(pio(F	����A�i� y�9��.:���ΟN{F�͎����3��ӆX���	�`�$�*x�にn��ޕ[��ȅS���ǰ4�{r�S�0���kI����vZ,�hlc�
�O�gb�xI
���N���^��;���\,1�a�3�%����q6B��繹�J]۬(���<��s�C?�d���
&c�hL:���jL�b%R���b�\��Z�G�r�����O��ٺ̗����|�'K���͇n�~�Oː}�����5��h��x
�8�Tx $Zrh^�`�{@��� p�}��PDH�1l����; �<H!�m���ܸ��
C��8w�cq<T��x�.$�X�	��֢��s���=e5���� �ڞ$���^�R+K	ҤyP�}cK�E�~�G�������Oʏ���s�tU0`��Q^z*�A2��V�Y�1���P8���^J�[�}��w�q���:u241����������Ͱw=�梶���#��;���j��������|��aK�k*f�y��՜���H'���:>��ǃ
C�J�������y���h�X��Z�6�Jcw�`qf~N޹��,��H��%���\�Y����*�L����!9��������>�+����a/P�����l���A�i]E�7�b$�N��.��'='s3:�`�hnK�ܔ<�ec�HC�����T��B~�s����Rg�)/�=�-���"���nm3�8�WC�V��ׂ���p��`��Z��zR��-��z�.�N�G�B@/�G�B�p�s�EG�=��~o�&px/њ��*��m{wwt�$��s:��'W��G�������䭏.�G7W���!��S}�E�t0"��ށ�"t�2>�ъ2��t�j�K�*a �"9��9r�-��Z,R�����h׷�{iqj:`���N?���஗��#����Z���0�b�ѩ+���VP�6���=�2��� +���(.--}����QN���(}�vX֛rksM���c?' :�dM�$�������#ZD��͵�puuU�i_���^���l��.$5�gE�db�YD��(Q��t�Xs�<AJ�ݴ<��si���S��<�&��7z�l�ƩRӒNx	�݄-��pj* C�ɱ�%y��I
�e�yU�e@̠��"@hг�q�u���
`��:�x�}�>�����
FY��}-_��TU���dfcE�����H�7�x �Qa�����&Bλ��V���JBi�%�,��Vk�@}��jT$�dH���Q8l�!)h3XN��SA�֋��~_A�R x��>M��bk�:��OXG�R�I��8o�Z�[��G��s��c��˯�)�|�Y�ڑ�>zh�%�����U�Za��4�l�wj�&�CB]�N{=7�ў�����SGB��;�;�p��ɽ6�	q�� qahm�������û����]�M���>U��̑���<�[o�E�4<�����mRS`H�d��x?�ڽB�����*�'��e��ι�K�W��^�O�}O�%��~�����=�~x�3H���ΓN�(��3��h�����!��YT���rX.�|h��8��$m�O�~D�_�$s�P��F4v9��qT5af�Y �`�< yt����'��}ߜ��g2�q��qq��u����Jf��iH���u��m�wY�1����v���d~� �-�S��ʅ�G���R�H��n���+%�^�V�\��6�9S���j]EmL�$���".�>�Ak҉�	�
Ѓ0�UFềoA�'3���}��%�A�5�, 5���%�'����d��^���Ǫ7J
r���~��"A^S߃�n�ƫZ��*�?��=shT*F��`7O��e�|��� ��%Oy�eX���T�x���=T�;�r��y��e�`펴�U���s�� Wo.WV��� ��9�d�T}���P�S��!�������yv�z�=��Q��bpGn]��^Qf��^����¨�3랶p(>��d�ڠ�ln7X^���_��Ym�]��.�F@@�i	���.�o�?�X�+�tB�������n�e�V�B	C?`!�z7?�A!:&#Y�ޓ�
��Kn��@\��c5��O��^�2�K�g�6Ҡ?��Ⱥ��8E3/ d����.�"�u� �KV��u�V�\��:h���|����h��T�6֥F|�}�\bN��� T�Gj�����*p�)�����n����H�m]DPX��:ɯ-��<{�}�q�Hmc��5|�û
��|T�@4������׋W���L˷�ޓ"��;YA���b��3J�;v�cx�P@�\�o���\I��h�9�>�NC�ja�ޗ_�3�K�ֻ��;_�����y�\�Y�'������⻏Gq���զ��|�*&Ľ+������N��"�\�η��JE�w~fZ�g��$�looq�x�q)�0޽qcz< ��{}����u�1|���σ�я� �����h�ϝ�yzy��)�����]I��V+ Pλ��O9"�W+]U�R��Qy�}�?��}�N>�ð�����|���������w�'�F[���[�m�W��n[�ڒ%՟�=zA���E��ai�N�^22F֢���ğY;q�u#w=��cM�#�9�>*w*�?�-kĿ Ey�{�k<D�
z��8����̔Гy�b��8��S�X� ���}�\�k��0R;{�lK�nP�!B輒p(�(n�UΫ~��9�ʼ�j�"�:t�SX�m���z���~���+��RQ�A��|�'�+���| �ޔ)�~�>�(����T��\�n*�X0��d�$u���9_k�fb�W'�++"E�X�;�m��u5�t�S�v�X!(���>Z���|eey0����-�j2($��ז�֥������Z��1�o+�l�ߞ�?�g!P���qCy4 b�˵�vgė���Fޅ�F6��J���H
REӛ�~z����)�jEE],9��S#�	��6�yn�Ѝ��[͞�Һd�G!籰�dhq`��a�uVٓ"��
E�%�Nb��B�J%�0�PDu�Z?'u>���Z���%h��=��� GN��}�f��_��9�L]HL ������ �l�j���/� +�r!y��q��>�J��B���[ι�}q�-Kt���vn6w��;�|�6���[�P&� �2,<�=���y
 ez@J?��@�dA"^ * ^� ��f�j:r��u�RP�+��3����E�"����)Q�3���*��L�Hf����r���nu�7ߕW޻DzO��y��]8�A�S���3(�u9>-������>C�{(������k��R�z�:ZŁ*�&I�j��u�'aO|�b�L��r��M����W�^m�[Nb$��Ó��
�^���y��4c;�n�����������!>q�}�L�$����G��J�&�ا9���h0"2@��:\�8?���>�w@���:d�Й�1���"Fj��̰���8���'�I�<_�y�#���l^�v.�9�2������<����\�R���Z �����] �䷅���,��`?�q�d���/��P���8.�>=W>������ex!����	p������[��5b�4�o�!����\2��7#[K�E�����DH���vD:�+|�8;��g*

���9P���������܅��� ���W�k�㋏��'.�����ߒn���4-)"t�D�y�B���<�8@i�
~�.����dg-G3��@�o�ѳ:�>a:�<;��߿�)�++Rj�蚈~S	�_�#�]��]�IO=X�w���ȔX���ͻ��w��0/?��˲��'�\E�<�������LI˂D�pmGѰ(�zJ�2(Teu�!o|���>q򿛩F��)L&6��n����\ �^�*�y��*����D�(�_ͅl2��Q`*3#<%C�����`�'�����Q��C�'6�m�h�qc!ף�t}���Sk�^҅<��E��)��2|�G�/� ���rw�lݾ%�
�f����J�U��80�l���0#�@H�&(b�4��B��EZ�]�Da��}��m^�`ъсe�R'X��r�,;a�<T�H���+�I�͖�GsCs<�t�ӃL\ah4 </��SF @3t� ��� �#KP�
���y�zF؍�:���9jr5���g���_�r^��V�6�D��gd�/��'����������,l����"���6ƪ��gh��.D�P�u��r��ս�6�9J������)<>�g1���u� /���+[aK�����)�766�֭U��ܔޱc�X~m��c�3��l��� i2���.�M"�U�K3�� �a�}/�b����&��>��н��}�ł�^�E�����:�Z�����켼���?��5�=�,]׹�҂d_��g�\��9�œP�HX�Ӗ�!̅�H�iv���i�h{ �tz������'e��Sz���]94U��|�K�A\��Q��U}��!F�9�%�n�~l�/N���D�8F�����|t����O�@x�P!=U����u�� V����yC���.wQ��N�;k��S����m��g�i ��Nz�a,ϵǋ/�1���@��[��������"���4y/,��qu1g���jxZ�|�)8/(����t������Eڕ�Z]^<s\YY���ܒ���/����NՍk�u��E�n�N�g[�b=��C� �.nh$
����S�2r��cչ���nW.o���L]�{��j��Z"�!���+�����7�m)�9߾rEAb�|í����uH�NC�^��9&�յ�:�9�ң� S<f�K!W���^�Co��_|��'�O��WI��c|�a�2'F���X�%��������z�/��*u�f�4��M+z �O�V�)7����.�_1�$>K��=��)Xrt��9��u<lk�GQ�	p* ��ZE)ZJgG��?��Y��������͝uY����ʌE���nq�6U0 �A�.X�3�|����)��LT����ſ�g 24_�����Q.X_Mp��2ɿ�M�]\��8��a�z0�Qh��z�J/�g�r���S�E.C��"2���2�^�؊ox^'P��������g�s�y��$za���$��t��C���?�
^+��w^�E�ۤ�Q+
���J�ݯ~Q�y�1��[���ߥ[��8#[��4�'��qv%�O� ��Ϭc_���L�f�����������D+� Gۻ@��o�h5c�F���Cw��ׯ�[��C���r���� �Α��3q����M2���\�"� eV�И˴�"��I����>w��� �����,X�=8�����^ӓ�� �� �� �����wt�qj,�=������k䥕+%2j6�jH����ܸ�IGBW�ƙӏ���{ߖK[ruOm������N������3�5����p��5�y��pn3ߡ'ю��i�#�E[�y�D=��� p4Jf|��nMCh9 �	*����=rHN>}Z�}�ʖ))D*�T��@�*�Zq��\;;{�Ԗc���5�~�3W��#�BA��W8-&�-,'a��d� VD�8��c>��=�	@c���~����Y8�o�)�%N��S�4A`��ǒC.#���r�G>6K����Q�gS�d6������W�6Bo�+�S�a|�i�����up}���2� ����J�R�[Y+�m����΂�c��r��G��S'�����O�+���#�)PA	ύ&� �Op�\���8���Rq�|.i�^ȴkΖ���s;�XA�KI6u^�|K�@J:g�����y�(%h�bP>ʅY> +JN:��~Wo�Nѱ��������Z��
���B·�����u��ũ�?��:w�������2�H�X<x�J�*^}�(?���ǯ�"�+3=q�x�Ӆ�{h���"�]䅊lv��'o�#k�4� ��{+�{q�-���"�������fO#���z�6��9�`{(샒�a]�&Jpq��i}�i�!��d_x�)����P�$��m]�M��H�|�fj$��5J��T��t��5�d[72�0f��#l�A�9�p`���Z�O.��8�,�7+k�����`��fAb����e���xk{���m�I�j��G���>Ba��Q�$�d��FymPY�|j`y��:�d�KG��
�����ߧ�S���K&��r]+����˙�c���y��_��e4m������\7�>��OsC7KvF�4NQj��w[pȒ�!���T�]�mn2<�0�yQ��)Ǐ�`8� 7���st�ْ�Y�il�Q9W�h���{̲ ���~@s ໗�p_g����~�$���E�ڏ���> l�y��s9ʥ�B�a�e���T�x�9�KeO�]5֗��d~aNnߺ)GF�~�1����5x�����XΣO���R+I��$����H7x���������C����J��FQ�SC��ֺ*�T��*��ŧ��g��ZY�[k�����l�-W!'�����n�	~L��e�d$zj'��wD�V$����ɣ�=[�p���!bD*37?ǯ8���W��� ���qy�A��b��.U�>1rn8o.�����E�0���9AW��wS���K�@�c���k�����A8�K���n0*<!kұT�>�d�c���Ɯ^c�Zӱ���6ewkSJ:�=-�����@~��۪�W��S}��>�Q|���Qs3%t� �5]��9ͩ2���?�\���ע���U�"ڶ���G���޵5) Rډe�^M*���R��!(�,g�OZ��(y��<�zz߻�NJ\03/���|�=���)��vZ�R�Լ��f=D3�ͅ���>�����(�	0��DIX[-�FU��>�ݔ��KE�����J �Pȹ��}IV��'�+��PV��.�?��o�g�.�N?��f_Ν{��
^ekw���lB�C�F$�L�p��
�QD�k��Q� ��ƛi[鿏����TF䨡x&o�`gjU�_o��)���c3��9}d^�P-�ݕ�r$s�������n��-I�r$�6�#�k����CvvnV�kSr���Б<n�L�U�s�Q
����J*�ЬF�������ׄ�10�zC+ ��vN��`{gü|�.Ǚϕh�`"л�?�1���K�B��(uB;+(����豊k`}-�h��'�\5���,�k�C���}Z߱3���N��g/˟���|��&ۍ��?$�^,-�A�C���<���M�˾��r'^�"�P�I��@b����R��W��Z|�0p���z횬�ޒ���t���l4�q��)�����.E#YR���?�z��u|�*��=L�_O�E��>���
=�6p�Y����ȏs�#p��U�����������ܴ�,̲�"*��lb/L�L����� E�	�~���р����ҳF'��BW��]���pl��I��n̼?��Cz��?{-Y��<{�|��'��9)��%ۗ�C���V��SAe$��P�9 1�Ą���`��I�0��"0�� �9��^<.oc�U@`�M&+�Cx8(���G�8M�먆V����m�\oB�{v�g�-��GY�ѷ���}:4��Q�u����W7�WmkP,`$��F:8~�=�VИ�.4����2}Ƹ�ڵB�$���Ha�)Dkۼ��
�� jˠ�����>�C�X���3��sg��W_�7�}_�t�k2��l���UźLv�-�cN"�{M�)U����O�#p\O ��sd�y:�+��t�G�0��k��]��v��Ҝ�����٩1S�

�Ǫ�R���h�Iv�r���:i��}�.���ʯ�_�����^E���v��k<���2@o�bN�G�y����ػszvN�mݢg�:U�ۍm���b��[�n����w��b��#�����:��V�N���9�����ƽo����^{On�R����h�	b��Q��jμUd�4	x*WD����C\$ ��抹ѻ�v.1bE'9��R�1��rN�p��<s�,N�u��ҕ>]�ʌ.��
*f-�ʖ���4�	�ѡu���Qr	�.���eac:Z�Q�@�d�L�u"'����Y��`�����c�ϓaU��A���B
�E�f�>���@�vw)�  *
à��ʰ&�gP`�I�l0\K���6u� ����^����`�y�)��'<��ܐ@̈́a7OE�& ��̢~�
���ߒ|uJ�9{\N�=&?{�u��k�ʭ�[圁�v��VP���N��MaFy!�7�{�_ɰ� ����3�`�'���}V���VK��&���lnm�M��ton2eJ$��G�I>�����d���q���A!�~�w�s?X<�s� ��σ����8�\����
r`8���2ljv�m�vt]���%��'g9��\������:f䧓�E��H��y8-��ϻ�ҙ�I��=_j���\P�vrnJ��������2[Q 0hHU�f�+P���2��V{̄��ˁ�����X����4�D��%� �@b˄] �S������#�����F���'�5�:�z8��0�UpE�'��P�D3W�`������aAFb�`��1sY��ad*0���C��}�3=��"2�o�~.?nl��Q�n x�u=�p<)��Zv�k�T���Eiw����cح����� �--��~�Cy���٬�P��p
zB�M���~j-˅��T�T��R�V�Ԥ�4#�^�1�������#>{tQ����ۻ��&$mYW���B]ά���^�N�>�����������E��`��?�V���G7��o�.7�ve'�}\�K���	K�2�Gh��>a���e/f�( DcD������RC*�܃jmZ�8y�n/��\U^�hM��_�7��Ϟ=%�J Y�-���$_���$�F�|�N �/]����~��{�S��n�(M�$��?�~�@�sCWB�.w�W�:/N����S	X�!�����B0/���}�=I#�f�ZA�-�o����krzi^^|✜=�$���jh0�/�,�{	�'4r���*n�(����Y*Uhy����ب\^�u��v�(^B�3�4���AQ@��}`|Rf5�����m�|ވ����U�ȳ`�Y�1�x#]B�
Lء�};��O�;�3�FD�U*՚�ˤ ME���3m�EXm8W�B$���j�Ka������q&fe��^�<b�W=?��!ti��˱�ˀV'�e�h�<M�b����	���zhQYO�4�ˬ
��K}�L�u[�Y ����3u� ^���l��.��ƎdG7ր!�`4`�c
�c��P�!6g��.�ƕ7�-p��z\�[`-�R�75+B84A�|Ҽ��EB��	��@X9�L+�:U�����c;���Z\��"�T��-��f~ψuLS̏�9h��W��3���e�aV��}�2�$x2��X�sl��C識�s;�;�����g�z<7�Ep�ϋ�w>ԛ�2BKVTw��� L�JQ*5��X P��XE�L��u��Gɭ[kR�}�gl���l�G�Ɩ��������9h*�%ꣷ���&��ʁ���Rw��YH��i!s�Rz7�����ZLm5,�X��pY��:�o���|��di�,]��M5�A��S��6q��{�X�d��y�z-�IDЗc����8r��'d�R�0���Z���4�9V�ҕ<�e��|���j�������1`�a꼨��,D�zI�3�1	z$��lnm�i03;Ù�C ����XckXG
���cԧG%r��f%��S�k�Z!P��0s�Q6�=P�`y/*u���T砫�|o�����8������ZB��6dHz�IL�g0�0�K!�>�Zm^�wG
��͞�Y�!�z]^�pB��o�/~~Z�����rs�,̝T}7���e-镳��ø6�l��֕�������s\�ё9�<�%�R���#��R��4��5䦞�k��<�&3*�O�:�QI�7�ڮ��ݻw����nK�n��R�:W=�l� �Q�-�9��kׂ����ˋ��߿�&���+|\E�y�Bg*l.脮6��G?�sy��9��g�J�=rZj��ˡ�ӈu�v���E������y�+�ޑ�7V�8�,�$�P���Rb�5�
8pճT�=x���{Ԇa�`�H�������^�f��6^b%��E��{���<~bY��ԣ2�77��`T]��ٙ��_ < �����D��
޼Z�� %�@��2��q�a�떅��؋ȑ�.�y��Լb��dT�Vph�B}n�?|u+��f�uGZ���K����#��r���~�)6�)z�P��i�n��}�g2���b����`�c.����.H��2�q`_A�+փ��.�O{' � �if$.;�&|�5�d�e� b_nD��1[7�:���{�C`:7W�BY�zkO����* OTr�w�%g��X~�����]��g�ᬷ(M��	e[[�:t�bن?��z���Ut?��g"��)H����	��|ؽk:�� 6��R5����}���Ar~V��:��݃88?��{�'A�<ic�a�O�fڟ?�����:�G��iXa���fa�X���G��Jh����u57?/{��67��N�Y�h�?��XT�B{<M��}���t8A��D�(��Y�oU�o�oH9P9w���&O�<"V���Ҳ<�:o�p��TM5&��5��P�� ]V�&���&��C�3������-�ih�f���7c�<wd}�$����9ܾZ�E_٢������yf��BJ�>:��lN@��y}���u�"�8�����D#B�!k'���y���l�X���'��N}�L�:PP���I�y|I*��l�����3���X����ͯ�K��zSpr�6������]y��i���=y뭫��Y'#
�o�Nc#�<�_��-�h���z�����R���HI��E8�?�d�"��<� �
h��*�Vx��f kR��ꕛ��p�|����E��i��G�,֥_N���1��FOu��� 	S��+V��j�|���,}��5}��SA;:���"�w(߱6q`s��┤,����V��kWeQ7��S���������&��P��k�v�+]�-�gQEU�%�=&}4�F�SB�M�n���{1[����Y����o >L��0K��,��U/gɸ�<1Lp;b�<��d@� �mE�<vnE�?sN�.-J)���>�(��l}^��fx6� \�5;g����9�-X,JO������D�N	�����؂��� �#L����xR֬�����~�x��G}v^ǆ����a����i�q$9
��U�:tH�
�0f�UT��T� ���]�m�t�U��Ա#\�t�dAb�h#8�0>�;��4���#D�$�H���z Ҝ#Ti����w��;37+5�}�8y5A*�K��W!��#�eayA~��_�Gw7�	J��@���l��C ���C'������:��f�zt�C|o��렃�}�Ѻ¢�
 ��ݤ� ���,�Ѐ�s�6=�f��NP>�Ƀ���8fs'Ab�3��Yz��p���{��ɿ���_`��9"G��U�ۯ���E�ա�^�*�<eYk�!G���H)�;����U����@ꋻ�����?��uhy�q��~�}���.���{���J��c��\����r�lP�������Ԃ:{B�Η�(�]�i������I��3UY4��-��F�oG
���y�G��K\���9B�D�M��Hx�|�����5�ix�������ۺNx>� ����5����=R����I�XgЁI�9Ӂ�x�
����8^ӑ�4.���ɀ�P�6gtvѰ�<� �(���cb�R�Q4�z!g�c���]P��#���:kmn��E�_���I��?���襟����Mե<3�{*��l�����Rw��w���u{M*+!��i���� ��F�� �� >�TI�^B'�]546��>�Z����MOeX+�</�VS�Ҭ�W�8�ט��i�5~�&�)�	���_8#��	iP�$�i27�%��[�E��V��7���U�U]�W�|G��o^#�-#�S��L�h��G�"�v�\��E+q��ВO��
W0�ЏY�s��x�B6����������{w6d�ɳ'�������omޒ�tQ�`uW@�0^�T�l�n+�H�C�**Z�0�1�0r���r|@7�7n������P��߰7����î:{ �1�H(.@J�= �����=S?Q�T�װN�*�Jw2	�7S�!@-��jN�&M�~v�$h�➝��1�	���:���Zˑ��e6��! �g0���FF�2\��s��{¿���O�Жy�.��l� �Ľ�-^�;�F\���M��廪0^~�=��կ���_��1�b4&�6J�=��M��=�E�E+��mI��;ndU���l�8��i��wE���T�5�Y�?򖬥V���]�#�����_�1I��<$�;G�يl&���9�`�������\|��/�㮋���T�V��ZB������ҕs1��Juײ/�\��:���_�W�w_����w9��r��NKj*Kx�ܕ|�!gO�o����Y>Dڳ����������5�	@h[�
�u� �6��`���c�"��؈k�g9w(��/�ߦnN�Xo�3�.��M��,צurO����) h,>:�\JϚw*�d����yL�$B�����:���%���f��RW��|��'[K�}l}~]Tx'�i�r]k�|�7[��C��T!ts.]�4<���s�X>D���-���J�ܕ��ߕ�_xJ����_���tP�HUȡ�ӛ�j���guU�}Jb��ζ�u;2�rD�jx����y�9�z]�;�8��d�57AD��{PE4�`�H���zm����7�|���E�L�'��.a�w�_)�<�P(��<_��r�("N�/L�Cq3!Ebgc���!��6��]�5{�R�2=/(V��xR0K�W�:��������,�0�Q����0\��,T[��K�ykSc�X�0l�_Ik����P���HM��rҔ�����xD�׋R
�����Ҝ��.KI=@��Rz��l��$q�a�uK��e7v	̐���3� ��a��o����B�b�]�m�&�� �[�"y�+�0:�+a^�IVS�X�;���)@>�W��Ȟ����r��-�	����
�`��! F��j�:|��L��3���ޖLMO���C "�l�S<yℜ:}���\���G��{ �����~��
#\�P�L�\� �	�{}� ��]��y677̂��D�M�Uu�=�>L�,V��ft�= �������V��r͖keZ�
���j^�?|�EyD��O_{K޹�.Mxj
y�������#/�0�����%�|����哱��a�9<��v�Q���~�Ul�T��ZaZ�ʜ��Ϗ�!��kk\+� ��u:��09�w���WJ-����d�nF�p�g�@%5��(��C�
{%�⃊W�����~���,��kf?wP�A�w���5��?������s�yٻ�Gq�'���~�T�ť�uyɳ�i�����k��k	w
f�B������L�G`�
�L����s��~�!�=���)防�sX^�X
0�����Q�����ܣ����E9��LYH�������z�A��V���{�R:F�V�����T�/rFz��E��?��0�Ge���6� ���K��u&��6T�@^�X�:�������]_�}��/EQ$t�<��iB�,V�=�u�� @���u��)��m6�������3�m�t�-�C�H�`X�8w��9��C!�Rm� +t�@ĉ��b���T�T!D���Œ��;��'��R���b�O����=��D8�zD#�O�R��oV8F����W\�g�����������R�����������_��b�;=] ̪+���͢�x�]���4�շ�w��i5�+i��iYm�@S���$SG1�p�����5F��GR���4Ŏk�-�㣆LIPA��y��zk!s��^!P�Q�9� �Ͼ�MO���~�(�G-���_��#�d#	,lAc��X4y�)�Y3LtE�Aa��~7v@16��FC��>�	��dK0
7�g����x(��
�֠��|�)Ϟ?%�k�K9V@�� ���sgӨ*��T��r�~{w���w�����8��=�p��(����\."��u!�>�����"��}��^���}��~@�kׯ������l���'���稂�`w�>͍*�P �\���3���c��-Z@�[���(��Ǝ���`�������;=,//�#�<B�o#�
��
p��o̒��̥�������0j����+m�cB��pf����%�IW�sD����3E[H}�H򞛞��n[��A��#/�9)�W��_~Y~���*8�Se˜�.�f#�$���z�G��k�/h�Hs�)��n��SOI2;+�^�
�5�x��8�gΨ0\���w�>��xr��	�#���k�9;�6��C�Y=�v�l8;��l�Qt���7~�cH �9y��'J�l�1߀�N����ۥ��=�ˢ���խ��E�v3�Nd؝%M�!�?Ñ�������e�9؇98^5��ǌ�_�%�NS�>$��_��ٚ�ΓC��~��l�d�8��Okl�P���<�(g��!��>r2����0�7<�b��(� f�,X� 2���'#H�I�qRz�C睄lgzY`)RUp&	��D��0&>x�}���( ;��Yw�bֱ�Q��/</��?O0�n0��KK����=�����J��	=�}�9��3��t#�@(\���P<�wE�6�0��qnx���`zPlU�����B��|� ���ɑ�)����uZGQ����((����}�z_��կ�K���~!���N��Ƌ�o~~If7e��:���޼�~O�V�JX�+�T��F,ۥ7�!�4t�6K� u^�q]��O�1��e�OZ�?�v�bd�ڔ��V���և�d��
�Q��$�KP����6�<9��Xp�3�U�zJ^�����/�{i3�=��x�Z��$�AT��o�Z��B�`��9 �Cc	�����VE�i�,��Q� �<�d�G�քc�h=��*�|oO�y�Q����(q�!�U�YX���9�����]$�[쫋
\q޼!IJ�����o���悉����X�H,g�g<����*b��X#�Z�w9�P��{�7��o�[y��w��Ǘ�2m��7��Y��x�?����;|d�ku[�	HW�*7���q�F1Mh�\܉-t�jŮ�F�� (Y5�ٔ����ի� �?�y��y���|�qy��Ǥ>�B>Ix?���9ڄ�kEꆯ���5Q,N�,��:*�N�w�I-�8B�9%jI�z�k��9%�9}�]G���*�JI~�KO����_�!��=ie*���\=�x��H�z2�,ġ��<iOqG��JIL�8"ٮZ�X3s����s���0�k(�rْ��v�� �{��U����ˍ%�O��g� ������o����,�d�y�K�_��kܛ���alՎ��i�A-RݟtE�(��`e�v}� ��^�������{H����|���+�����b�Q�VU��پ-%UGg��O]�������i)���Z��A��n���F}���dD��3�A]j��Φ�1C�<L]4r��J���>"bT0 �춒�\�&Z�vo�3�&g�e�J����/_�m��ɂ��������������a1b���&tuµ��^�`�[Dz���Z�����b�4��G����P��O F��V���c�daq���H����0����=�ϣ�F .y�E�����2E��[U�//� �U��qzFstz�"��ĭPd� �F���;S�2Wq0��&�݉�����f�d��$�LG�y����g�˴��Ko�I*���]��dk�+Փ�KZ�-׮�wZlԱ�@sO�S導^Tx��.C:��omg���n FQN�j7E���,1��sVc�匦'Y`yy�T(���'��G�ŵ�/�iv-�G�i,����̀�ǌ z%:�Ub����ִz�-E��Ih�B�tg19��~y��q��>��44T��f8�b4���{� �5J��
Zfs�@�������Eټ���պ\V �W�X�q���ځ���� �}#]�/�F	����YLMT��%d�������A8�*m�r��aZfX/��3�Ex���C��O���E{& ���_B��Z��7����So��x�����+{����B��T�Nz��mz,�uC�7m�v���`"��U,D�7]x��&2�Ĝ~$��ކ
�?���V�R�}^Z��/�a$�Ν������C�,�vaΐ����4��:�`"�Jv2�Lc�a
e���ܺ�Ͱ[�X�y�KuzF��:ha�
��!�Ɔ���<�����[���#��	��n���U]4YR3w��������g=Xqka��n�qMF/�\^8,'N���sO@�XQ�����!�nG^T���oܐy����q=����h��Z�8 ���Z�^����`�@�������:C�[w��d��R�<���>���o2l=vo.<q ��(�+1ǩ�FC�i��NWn��Ji��e�ۓz C����8	�� �Ľ��ğ'+��~L%�Q�8���?��S�;/�樑xT<��&�@��@�b)��*{=zX�r�I�+�es����-���^��Q��t���������Ę.�rA8��L�����s�s
�А�%J�=O�1z* ��"�ǈ��Pn���*(��`�[��?��W��qpC��;�G���A�#���tׅ�}R ?��$�}���+��P�x
l� <��[����s�K�(��c�+��gϞ�.P��NO���eii����'�m��~o��Q�74v��/!;�1�uǣ�R`�]t阋U�y�C*��[g�{�=�,�wx��BJ�$�Ǹ�P#ɜ#�Q��7t��4d�����#������+o����ĭ�"YSGW�ޓ��_��ӵ�N���=�Y}����"���5g�u#k]��8	��� ��r:"�K]���Z�:�H����(��~��_ٰ3���g�/�M��B�#Q����Zv�"]q!���`tfDv����s�]�Y�}ϤJ� � �;H���E����F�H"T�Z�Ҳ$�zo��b�!��� ��Ȣ�R����řeZbK��l��T����AGT�
��C��_�(���4GC����>"���
ΰ1��  �ǱA�7�)�W�R+
�#r7P��=��z��_ˏ~��a��6!65����>���S�W��G�!γ�qvv���� z�&����h�<��兄f$��:�Q�9>�ŹyY��.�t�
$������ث�W]շ�\A��VVV8$�O)H� Anʫ7_�W^y�B��?+GV�y���(Νc�%@��+���p����]8&�"��oZq&�6��:�aU&�*?��1��2�r���o����r���*"Tu���+ץ1X�/����,-����˥�dzꐴ���u�]�A����38mFG@ŘQ�n#���0�����B�=��n6��X�ͻ[Rjt��#=����܃H��o��6�GO�:�����ArK&�\�}�S�|ŁE[�NAޛ��)�Av��o�5��.��8:������{���f�W<���L��;�Oм�z��`��/|H0M$�g��3�[���"}�w��'��i7�n��.F�OTi�*7�ޕ������y�í��(�L��>�>gǑ:9F771����=�'@��v�ս>E*���yU8U i���1�1R�-�%��]Հ�ۑ�
�KO?%!x�ЕJ?���#E��u5
��,��'�<4TV���t��^D1���jY��$�����0��?%5JY�ó�j+a�4�����> 8m���В�7�	\����"�3����"�޻$7o�T|����k��#�Q� �b>��A��5j7�<�� 3�Y�

�*r��	Wx���|ffVf��C��>��V�������I>���p���B�k׮�������SvN��:v�=����w"ٹ,?���xJ�$z6-�2��s��#�"P8��{�*tt���N��<O�|�<墵P�S�%$/��ZG��rU�J�:�"7n���K���S���@��ko)Kk��Fء��
Kr��k2�k+��uy�'-��ڹc25?-�;���B�
ۊE�c]��cd�,>%Z�ׁ�ܢ�0�=u�w;���nۓί�́�t(0Ti��G��2ꐓ=�@�yh
��蓤�lgd���	�6�^wy��^���gŭ���Q%�g>F�H�Q��%NX���ߧ��T@<}�� Ÿ!w�]��z]�?&��i��!�B�ͻ�<�I���ƉKMٳ]�q,?$��/䭲�:�,��\_���)a��ȑ#��0p�+������?՟����5ZGXȰ��?9,Il�NlU�h_��M+(���۲��m��u����q��!aad�;kk��2vI̞Dc �{��ꃇ�8���L]n�E��ba䁂 ��1�(���+PT����Q ϝ?>�芼��[�o�Ϳ�
l���oʷ��myA���O]$��
4{m���^����Uq�v0Ok9�� FB�*<q�ay4v G~	�K<�9�m��ݸHF^_�*G��?��ߔ?����I�4�G���r�#��'1�	��Uc�ܮw�����(ϵ�5SQ>��צ^=z�M�B!��/�^�HM�\�p^J�ΰ&@�yk����g�V�Y<�/� b� ���'�V�������*�-wk��|Ι��xH���Cz�9ʒUg�}�0�{�fK�i�~#e�Q}�jQ>����
�@���Ep9U2�j]._���c��pP8���Pq��$p�/�{~��	�`  �Ϯ����R !`��<�B�|���V�Kg뎂�T~��_����W%� v�TA_RS�5��xZ����~����F����S��[���N��o�
�r~��P�8ر$L��3A9���~���C���jE�UX�.�'o��[y��7�������W��E��ٳ��pX���df��!�#�(�:#�������2 z���S�N*-0�iee�� �3sK#�(s���m9O�K�o�9p�*uM8l�y���)o���|�{ߣ� 9�'��������ɓ.�����o9�=4v'��p�s��^L�0��2M8�n���p�<��9���@���4Z�|��V��'�粡��F��x"��9�hM�߹E|Q�Q��v��5��ʌ�I޿��������F�eL��l�,� ,HT*+��A�~ݾn�.
h1N0{�>{%tb���#K��R�mG�	�	�o����C�_q�a�O�<]���n��Ń-���G��db8!L$��.��v���)����GO����3��Bc��̪�?}�8{�������J�%=��e�p�r9�6Ii<.	��FrE�������=i!�����ܼ��K�ӟ�D~���o���u�B%�	*j}e+{ѧչ�c�%���Vo
aF��sV�;kt�W��+A�,��aQ�Io�b[9�������9p>�,���-G�-��f�H�j@�B
?������͝�-*��@(�
ll������o������D������� �K�H/���@������L���+�L����U>?��]��'�;�F�8v�9[P��W/ɑcG���G��zI^�tMv�}����y{l��ꉺ���Njia:Z��G��Vb��LU�ë0U�����¹u��0�3��{�3���ޥ���7�!/|iJv�;���+�w79�
���[�A�$���p\j�e*|���>�{kL�0N��^���~�����j�|���W�w�w�<���y��<�y0��'������U=����9��8t�#]�V�}����L�
�²�{�� ����e������P�c�d���3�F;ܮ������R��l�!�p[$�\�Ň���V�uB��+�?+�?����[���;�n#���G�
z�U��0C� �P�9�2^x� �Ǌщb(`T���tF�C BYG8]��}��&D��znD�`����3b��˿��~�����y�w�k��A�<� dp��o�k��_��v������ yہ��bьN�)��@`��/���_U�ryy�Q���Ü'D��ni{>QP�`9�3�H��[�Q����p�"xC�5�@0�X�����'��c��s�='/���S�����ߧd�@���j�*yGp>��ov��2�T�4����� ��v>-���9��-�Z���5q�ܾ!����]�w?���^�&E�э�=��t���6��k_ ���I��5�>z���IO�������ߝ����@n�Lg^n�:�a-�]���B�=j�)�����g}����k�=�Dƒ�<�y֊��0��	T�`��L�V��������<]`�-Gm�>و<�,M��,_*���G�� ���#_��s����tv��Ǝ[Z���C�H�;�:��9�X����1�Bx��J�R����l�~{"���B��0�#�Jt3��P������/&?Q��vY�e���{h��V����A����h ;b���5vI��N��[�l9ʱ��4x�>6������Z��nݒ��n�}l�������A� � t�P��Y����Eu �c�}�� ��6b��<� 8�J�����������o~����O�t�F�0~f�2�1�x�|Yxb|�[X7u�C)C�#s����t��T����R$ۛkR�������0}��d��>�yi&�˒HI��;M�R�/�
�f�q���k<�AG�u��Xf"=�����s�ޱ6��YB(���W��_��<����F��]����8y���^Ā��XgL w��w�Ȃ�,��V���G��ދB'�YO�=�|q��~r��:�rf����w��*���'+���1�|������HF$��g�J�/�/+G�P��t��������=A��Ύũ�*G�-��A2E*၀М�<��0���5J�x���H\�{'�3D�1TUy7{U��O�y�<w����C۵ASz-:�:q�r`ш�c�� ?�1�~ET��"BR�I<9��w���!���$ ����P�^S�S��,�r��=����~񲂥�3�c}K�kt}�N�%�3.C��,�X� sx�=�:�F��w8�Np^�������s�=�$��Z
�)Q/,��sp�`ض�,��3���chxz~�r׆����.�eŋ��:3<�r.�o	�	����]������S���|�e�Z"�.�Y�鎐���/�+���!rG�AV0X���
m�N���P`���c����ڭU�X�*a�&����=Yy���o^#�`�kf��Q�J����&��ܑ�{F�4\�؟���'0*���k�BL �mmqͣs|t����;)�ٲEm�9p�7��k��,�n�ML�֔q�X��`Tz�ȗ��*��`e1��*)1�ج){C��ˡI�v�^�}�+�N�W�N�3a�d�Qd?]&�@�IM�_B1HҒ���g�KO�����ͫrQ-ʧ�~�׈уX���&灑�a���z\x��V_H�i�l�|K<������������.-��	�޵��Q����X~�V��ѿ�Ū�[�̥��uB�G��7�p���{��[��C���r޴-�����T@�#���<Pt�o�Ȝn̙�y 5���@P��!�V5w���?'O�4��~ `wbZw����:_� ���TO�gyiIju��t���l�z_<�z�z�3ӳ.?.�7�~K~��/e~qA�y�i��,�����
N����ԹA�]� n�������m�$�['9��м�3*�����F�.��|?��w�?)����ܔûz����7G�ˢ��O~){�S��k-p�`�4�4n�X�1/#����gaIPT#`SEҚln�J{箮�
=I�)7n�xe��ޭ�r��(�鉶�������~�k)��C�#7��K��+D���~�HH[��w}SCWiF�y�O7��B���H��$�c��hw��X���}a��Yo��퀰��5��a�k�;�=����ނ5{�I��I�h
�r�h�g>3�f�V�;1L�O�*�-A��X3^���ڙ3�U��_�$Ǐc�g�����g]#��V#��;����a�k��b�[���F�;Ó*o�&��\È�rtx�URX�*�監ר�v�º�%U���#�
<,*_n|(����g� G�u^��b=��[NG�,��l]x�M����uV8��/�yta��H����lӊ�s���U�Q�`nЋݝ����H�)XY���z��_��~�3��K/�zfyyٜ
zߋ�+�r�7���`�Ix%7U�ó���#׏\�æ�l�12c]e<RO �N�z�E��H�@12R�P] 9��x�;kw��_�U�N���ô�_c�w֭Kp���B-)0Z_�M=��E;"]hFA9�s����^�Z�S��������?��xϟ?'G���>�l��������^B�L�� �`vs��,N�FN����b�ox����Z���Ԁy���a�b�)i���v���P��O��5��C����D�N{Sj�gE����B!�z��V�����Ǚ�9i�Z���c� :1ND�����S2䜤�a0��P��3�`-,��64ʝ���n��ӳ�	E}���b�R���ze���ml��$ ? #�1|(�7��"�sN�H�Aؼ?ir$u��$pLGM�L;���jK%�k!䧨�w�~L~�s�}㲴����味�e�m�m��`� ��z'�	A�&��C	=���xn�wY�\	<X$�T�R��4��cS������W�J���C����Ӫ�69��� �	ϙ�a�Ce�sc��^�Ώ���M�J݃] 7xA�� |�7��S�RPy���^?P)P�de4����yO�<A!r��n���%
�P�+H�(y"����L}�
zt���w�L��=�T��v�AXe9�W��g���S�ƿT�
��ԓOʹ�������7�Q��s�����Hѭ�g�Y�������B`���Kެt���Bɤ��d�(*��ܖn'���{� �����5��=�r�}��z�ށFHf�2��h�6Br胬Q�x4�A��Ō,K��y�,���X�"b1t��KU׾eVU���}~�yߛYHaG�|�KՕy�����=�9�<�9�]ܫ��?����wl���-��C�7j��+/�Bj�	$|;%2��W�ʅ��ӿ��)�'��"@@������^;��}��]���]v�YV�7���ۍ��2�\�g�=Uf��E3;v�b"�f�^�"���$|�����[QL�?������y��o���B.o�̡&F����k/�fۓyv�
)x�����z7fo�%�t�HtC�y�"�y˱c����П|PA1����˚������t���f�>������Y�y�n��䗐�I4�t���C]��K�ϋ��Rſ�kTc+�Aጯ��t��������zo��\�����?�~��׿�Zkk���|]�E\�b�ؒ��ݓS~<�w�[� SHU�>PO��F��*w�ݡ�n���y�o����H~i�k�e���=1!���u�����`��/ ���yq��AP�G�����,2�+k����J*��l1�O�*TfgUa��c����N�g����2כg�?���J��
�%�Y�͸�?�b#�w_��*��K��ɇ@;
�R(/P���;T}��f\����K/)q��\�+�y���1%�^�n�O�g?�95�`���ַ�Q�U�o�^��r��i͖�i�u�*]Z�����K�i�b��ՏKS�:�i4*��Vs�8X�R5J�Wϝ�]�a{�#و��_���׆�2��*cu�w�]}�?�A������b��h��ρ�*:tO;�� ��b��B�֥ns1�yY.'�(�P�ʑ����eێ|�W�ԩS�9�$B���BY�0<�م(��:M�D@a���x�R���-�R� ��/��"��V�6��'i����u�0qw��K��K�ѵ
-x�8�Ss�;���M�z��ػۖ/���ƒ=t��6}p�@h��%�| N[��^dxڑ9�;�%�npcc���s�W��ىli��n�NM�(����fg/����~��}Ⱦ�FS&���=R�dl����Q���.("��Dn��B�zaL��L@,�(��It�����[Epr��^]�:툯ıDdF{J%�KɃ2�B�d�`�P0[ik%�>�(��|��]ᔕ�e���� ^���rq�8uZs���B����/��=?�o��������穙��[2l ,�{����� T���,p����U�z.w"�AI��d�����nIj�n0����+s���M��6R�ه>�9����g׸��Y^Öd8����XL7�&b�U܁u7ѩ\'f|x�F�'<�^�Z�(��imJ���L��E6��W������8X������/SI���kU͐�aF���AR�3�Ř�n�ۏ̳�F�#4��0����8�����w.����\�����$4R�g��M��7n�/����.���po��{7�����^W9cc}~8�\���k����v����*�zN�e����j}g1�Kր���^q�8x�>�я���GQ�Hcݖ1p���W�*�X��U|���<#V�X;��7r>iF)�=�x�3պ�g����H�����t[� gAӦ}�"`�=Y�9倛����yk,_����~�'���L�E ��|���u6�<�l�؞QcSK�(71ف�`RSPf�R9<m5��>��=-�����J���ܳ*Qn�����g�K�z>c����'�TU�9�Ϣ��>9�W@l�A RX�����ʪ|�����C�1�ea���$���X��Ӈ]�>��`qm3�} F�!�$B+*�f�.Ǜݥ,�D���c6��d6�D��a:���> �`*H�6J�<W��i@�d	��4qo9o�-�T����9������a�L)~���v��{�3���=�Ѓ��W���jҸ�ʎ�� ��� �۽aO��Df.��J5���bd�m�I���\��2ԭ�1��E;�~�N>��<|���{�V�`��7lueA�4���j��cWf���͸��K�.����@���l����,�R�f!�
�OhjhJz��LJ����@�;�r
.�u�~m	�Q
k1g��8H3c�ݾ v]������G_�����w�b�jI'Ң��#�Re�4�e�����;�ntb��d��l�o�[^�J{ّ=�:{�*�-����}V����U���X���^�@����%.�)���bv%�UE������7 *ˊ�e���i�{���|�=�̳��x�>:R�ب:���rT��CM^% �8i�Ikqw�KQ�	�y�nL�O$:�;Ν=�c;v\F�R�c�ez$p���D�-��x��3�ͻ�E��=�E��� >�L"7@�Tbϭ��&��\�a�Qy��3��K.�;��1t�GI����� ;���]\�g[J�(r�0��?��?��~�/������ox����n`!��ӬVW��zo*�/�2c��2Ė$_����������3)�QhQ�4 �!���q7ڵQ���b��������M����/mn���UM�Fq!
ץ����v~�%���'������\���iT.{��q���D�&��C��k��*���~b�������?��v�����c�ʗ�l/>�X��w:[⨒��N�7�q0���*��R]	��0���������=�v�7�~IGۉF����B����{��F`�K\�<z1�u�\�$(�q�q��^.��_}�����7{���=���{��
S��3d=j{ u������N|�R4�)С�vS3P_���,E���R������m��B�P!�._Aɇ�1�復єo)�X���j{'F�����}��m|�X4I`�%w� iE��a?���J��[���Ep'�z&�ni
Ȧ�zo����*;'28�'UM:)���rId�f����?�����#{��E'bOܨ@��q~ضf:�w��tXQ�K��6t�c�cJ\�tI�;���i:��Sթ��Zs��#5�tl��.?�a}'ɋ��#0���uFF1x�M�����$����m��߃k���E���\B2}���u�7�}�ol��M��d-� ���\*F3B�&�n�χ?����h��{����P0�b!��l������$�$y���d�2�,�gxK�6g�,~:t4�N4xь��Q�C)Ȇo��:��ټ]��e�=|��'��_��-�}���d�6񒤂��'��q��l����NXӗ�Y~2������$���'$�Z!�Ԥ$ݤm��^����d�N_Cee� B�&
�W�R!����%si��V�F&&mtb����o�P�BQ�)7�,J#���ڎ�N������gYb:���BD���;�����}�+�;��[c�����vu� �Y,ͭ, Z֜�v��' ����B�^�-��g#��.�#榷:���fQ�t:���z��{WD\�ϐi�y�ư������V����VS
� #�щ�\�^�3j����ȊA*���VC��董B{��q����eCi�
�\ i%���G�#�u9zT 	0 ��&�Z��Xđ�w�����|0Zl2:��J̫���@i��ۻ_7*����\������d9��D��/�S$��0*B�#}H;�������t���O��ML�gFO�(c�!,���-S���I|.�Q�(b��ŘM��1�WK�p�m�0�*�2|}6���55>&���s��3fox�>��O۩�E��9h]�����<k!9u>���X҃)�a�E�&Szida��&g���U_;Kv��θ�7݉��ݻ���ф��|�����|�>�g����6�g���o��3S67w�.]��{L�2S�G6�b������d�Y�M�a�ݿ- L��=
i�y�����n�ث��J}Ǜ'�Q��oi.��H�����\��_)�������%�G1���]N�Aل��m�iDq� �wwL��!E�m��E���t%5�Ž����t��v7����-�׿J��� qs�r�E��d�O�<a�y�1ف�ss�6l���F�a�ͮU�l�6n��������VA��e]��1�.^�^��q154d�bK�uI�#�zp��j��i�S<�-H3�[��u@��9����a�&�Ui�������������|��T^�8Kt��6-����,�u̯e��w�RT�`k��C��N����n�_d�}'�w������߿�f͗K�8R�n�Jb��9�f��������}�=��Ӷ���r�>j	�E;J���%W��Cd9k�ʔ�#����zD�M����V��{HS�?T_��%��)��~���R�~�'0�!d���T���`/��������ʂ��S���{���!2�"�O�d�f%e��7��	���W�����c���&e5Q�!�&?5<(� ����ڞz���������׾���w����ga����p�)�ȞC�E���s�����iV�{ �A�����V2���(A���I'��� �~��[�6k��
��>�C���]]ZS�}hj�m��]v`�Ϩ����fgO=o{o�Ӫ�m�q�C���w�
�e{1U����e�J�RS�=Tb��=�ZP�ַb�^�n���Q̯^&�M"��z�@����i�_^���y�0U��Ek�,/I��$��b/6PQ���-����-�� �z��dȠ�=�|���=�=R�X�����ٻW��1Nt�ia�BllE���J:��	�v~ge�NXJ����萱��������������,/�yJ��b]H%�h���Y����Q⛞��s��Me@��.=^,z��ܭ���P#pJw��B���؜?_^^�q(9��)�B�<q|��i��IW��� ,6s;�0�S�|΃������3�qƿ#sH
it@����dJ�T��r,I!�Y�߭-���� r�	�����R 1ZiB��I\"��#cы�.V��.R��Ȳ�+Ѥ�si�ı�7�N�C1͟�@Mc��n�m�r��{�ٛ_g����ܠ��3�S:q���)&騎�q�%�B/�.(ٶ��HI��	}L�'}},�㔫�v���xᢺ�z�AhV:g���,p��h/}�K_���ۿ�����W����N.�(;ר���J���ܠ���e��� ���� ���p����!Ӹ��_�=24�⊺�;���;��(�����s3v�Xǅ~����*@95�u;�d��C���!>�g���[�g!B���R>|�1��]@�:�k/E����v��J�\�T�:Љ�S�s�i�cϑi�ϗDi����D���E������ ���5�D('�<�U��v���[n�+�.���9�3�˚�N�h��i����= rG2���K�Mp �h��7u���tS+w`�9K�;� K	`�Ğ��9N�Z��Ū��8Z Œa�R�O���j������y�q;w�~�@4x�4��/,:�����0j�l��[�^o�2�܄�5�D�wf��+u��W杆��H4{zz�v98��K�+��7��O�������H�1� ������n��z/��m'�ۘ�M�����M�h��=<�l�TJ�Pg4k�c��%`��e)�{�y���x e�Z�"�W ������C�"3�m@ڌ�&h%0���g��Fku4I�]���:��+�d�&�P�km�2'���S�!"�k~~K���/�W��{��~@ vpw]`\�Z%@^n�TЙ��BpP��m��h �	����|N�kb�@��~�D�qb��`k^�f�_z���A[z������{н��G������ʅ�'/��]6��x咍S9������(�1�ݘD�?*A���1A/����ןb�;�Њ�|�b��hY��޹�o�����WhZܘB�#���zj��H� �A33=��x�Z�!���h��Z��^���ݸ�g^Š���cT'������������h4��lTi��Ԓn�±��	���);to֕۷w_d�������o�Ư�׿�u��Y���=*+�O���˂��v�7Y]�)~,e��=�2�ǏO��|E�jE�eyI�:��0�����1'�N)�+�(���b��p�@�%f�,���v�Ã3�L�yq����2(���D�333��ϝ{�3 [�X��/(�Y�$K���'���y?���%������D�7���G	g0M��z��K���-o�׼��v��a��R����p�)(�9'��9�۲B*������ L�i6�"՗�:��lʸiú����UF��u�z�JC��;���#��@�� #MmA"��+��S;[���U�#���D� dj�n�7u�G�刚�Z뾐�lcu3:$wM�K/<�)�}��m[8-�,���m���
[�}{��Ye�閾�e/�C�ح�B�\���hKƞ�uD��7:��u�j�s��݊��j;�໶�Nn����U�����oD������^���#9x��-f���μP�QIA%�R4�Q.幸Y+q�l��f;�i�
"|1�_[vu�Z8�R���C�j�Rd��k�}`D��(��A-W�����U���,%�]V�Ξc͓E�����m�,��_��lnnNt����&��@����9!����Ƕԭ���;:?��~;��=1�lK
`b�{w���O_.'=�N6�$V�lkw�������9K�a�����jK���ѱL٪��D�lbl���^g/��Vko�+q@�`m��z���_+�р"�E�SN%��ܬmNm���:��Q�~k�?K�d�kS������s����o��}�c�,��޽:��?k��"�R7�Ԣ�/ʺؿA�85���;�ܢQ7��(kH�͚���SPŲ� "|����2���H0 �Hp�)d�!u�^�A6��T�H����7>ixx������cirH�#���m���u ڲ��s�v�7*u���bԊn�*){[�1��T4�%*eܳ}�C��ߴx��������IT�X�^|8�&���tکrU��U3��{֧��Mm�[y�Eb>�X�߶ �~�^z�v�_�������<e��܋n�G�M�JcCM�C�Ah��^�f#�<�Ac��B��-E�Y2��T�	ٔ��B�Z�\ś_�]���,t����śa{�U�{���Z��b����N*�5�WI�,� ��Dq���+���o��#��J#��kZݍ��<�j{�mG��q��/��ġ���){����B�?��ܙIT�!u��cK9�ݿ��Z� ,t�D�OYlX�$T�^�7�M��8&�ڹ��u,��}��!��ɔ��g�yV��p�~�Q,�����6����΂���`�}��t w�v���	������u���(ו��,��|�{�g�s>͘Υ�|�0RD� ��yߖ@h8s�y�!����ܹoL�Q)�f�vpo�9לy5���Ox����g�iϾ�Y���{�&4<�ĠR����&T�!J�l���բ���@F60���æ��537�/�#�#�܈�����#v��I{�٧�������}��P_�f)�v� �qL�1eN�0T��&����Cw;W�T��d��/�S&Ck��wh�{lt�jw�{�]�h���s��Qw��裏j==����S'_��zH:�pM�L���h�S�Z�pFY;d�0�#�g�<b�w #��h
��m��2�=ُ���ّ��p�!��+;:�lXd�c�T�@��@�{�sD"��֞2�

j�2�1�"OO�[�L@$^��Ϝ�OQv�ۑ� ��{?g��� /*tn�f��>�Z�@����$�J�$��j?X�3���zC����{�9W�\���<Y��'���ܙS6�ϴDi�nW`���V�$��X���������C�p�ի֍��ۑ���騹�;|�������A_=	Kg`��9G�Z�ٶ?�����z�-��X[���f���o�~��u���]ֶ��t��-�ow���4t ��++�����~В2�ijJ>/efl;�)S��;e�20?�_x����X�����f�z���
���O�r�Ft���Ǧ*sف�[�%��:&�S�1]��a�w��'���眳���]lj���L�Oa�aG9'�������P������lbT���FK�.=@e����s�-��{1^��N~��?/hB��ch�J<�h�K
 ;i��/�`�K�^=�ԓ����ňY�_TE��9�w��`��Zݘ�r:�{U�R(	�lgv�Şc _O���>�=��'lk�=�����l�g���:�ݢ����;�_���T��s�_X������!KM��;,�/�����l7@�8�sM�C��ɛ��w��XW��&t��x�Lk{")�V�j�ʰ-9r�XM\�������X$��ŬN�b��Po�ێL��`g�ciwg�a�7�TuȊ�6���w=�=t�1[�;k#��9��v�9�P7N,�Ņee����
zP���s��dʩ���c.�d,�)K�0���g����گ��=��"��}�$;$-C3E"��������h�N����<xX3�=2\�:�Q�?{�\����1/���iS���7$\��(kP�Z�6�m!�M�v��Ȧ�z�/y�g��EWK<�ᑐ`p�BIaځ��s���煑yٝw�߈y��� �ll�*C�n��.e����gϜ���y.)�˛9�q ��|��U:\������W��ػ�e�<��(��=��Pr���W��݊�"�4>*@�~�<V�jw��{SU&��n�ޖ�j��l����n��.9��������kt�>���iD�P}�m��Y�u�E�K��k���\��u_�5Q]���6X-��2F[��F�'\�8�������j�ܕK�[/{�}�{����A��sg����K"_:e������OH��رc�@btظ�('`G�os}�����q��0��RS�B��4Ƣ,�F�NG��\ܞ���!0!C��Iu9�,d<A�T�3b�R�PcV��+j�j�m�*#C��kXZ����j�h���� ���g���ު�?��8t�V.х��vT^J�j�Al+���Z|�u-��p�J�����|.:>Sٹ��4P����\�TSH�/;��e�r��h$|�������ܹPG�5M�>MO��5���ć���ﳡ��//�s=�`��k��{�miqH�;������-w&������ж�GWTyQ��R�?'z!p-7P(�Kd����4-�H۷6m��~g��v`���ݏّ�m}u����6Vc��X|�ueW6mrj,�@/�@�~t�1��N?2��ѭ%�x� W#� Y����	RP(W��5���`�_��د�����%�����?���T(6Р���u��{��E��M%d5^�$0�e��|!��j�{ت$���d���~f��ەA����E�N(9d9�[Є��z��d)+�B�����ГPޘٳWA���H��FF���=�o��nn$T	9�+δ&�:���nvi�Ѓe�+T���v�p�ڔ�xm���-�\Z�� �G����ӧ�ڙ3���x�>xP�53��XԴ:dҬ�>ۍ��_�J���v��x�zo���/�$�tkt�uK�vpf�-�-j\�k�G��/�z�
���>����6��Yk�6ljx�Vg�Y�Q���!ߣ߻4�4%����t�#{��������)Ee���C�Rh���,?�gffv=����
7��C��4��u�bt�I'[t��*yyп�V1�{� ��mkH���A*�M�^�mgW����b���3���ڰG�:f/�7m�V�w��~���-b2�g6�F�����C��B� �!�e��I ��Tm�t-لR�l��y�����=��O|B��y�+�ڴ,^۰��e(�ȣ�0* ���b�\2W/WdA�ܒ���)���F�ű '�?,F���I�6�Z�Z)K?��s~|���%FIٿ���fEZ���0{3(���{�pRN�����!��s�m7��$����{V�r��0��K�=A����[�}�O���Z�t��٢2��J��cA�'��;��>�<�r��g����7ُ����}�E�����J٠�ݝe�b���A�Q�[�Fsc݆|��G�dx�όڛ��m��O|�^u�+lme�>��/9p^�Be��n���������n����R6�9�y��~�up�ү�	 GV��%.�m�U0�V�4$���%���S;uꌯ��@�Ŀo�;w�ߧY��W�f�}�.���ʳ˥� �E���[][�Z���'��iIP"`U�}�Iԃ�5c� ���^E�����WT.'M���=�
 �~�y��t� ) SՃ�]��$^�:V��σ�̟�\X����3<k:o{�^���}UK��,s�JQ]��|gUZt�M95"v����[d"ݑJ� �$�U�����T�ZL�Nd!9>`+?��k��h6��c�N5x�9{���ZP��{փ?N�WG�P�4��<��"�d�`u��ON﵋�gڍu���&��4Z6Ps@��Mw��{��ǎ�:ih����cB:�W�R*�~|�$Ս�ڼݺw����G���_Os݆nų�(�N�6T7���53����m}�lh�qt1k�u;I�?��,���w� �v�\�\^��p�#��*Ф��Ϝ��#�������AO�T�c?I`{���k'��$�&��g��P2����:����)�`$l) ,@�}���6�-�e���.�r�9����l;�^⯸v�ѻ��*j�V��9�M�Z����b�sW�9����_�/U"i3���"|J�Z�Ɏc��;'N��_�L�Ã�c<O�}'5H\f�����2�) �����o����?�#��7�E�4�\��V�<)3���2��8��a?6�3q�>ah��"�ģ�L�451jC��-5�<���m����|�m�{��*��?wɖ$�6|�ϝ<i��C�/$�ZH�@�	|(�U�6"2שq�A	;�9#|�gߖ���h�Z�?�"۶F7ci�˴�XUY"79��7�8��R)VC&�(%k��M#�������aw;lw�g��]�C{���n�ZLL�X�XK���6�@k�������Ϭ�]�OI@�0��Ҭח� ��&�w��1~���?�qw� �=�DIC_h]�}@�">��&}�"��H�fpdp@�&�esl�g����`VY��ߏ�,��?t���3n�fgg���"�"���9U��t?�}���ͳ߁Y�<�)��0 ���瞓���pJ�$1n,�<�A�d*��KR*A��8�̳����H>2����,����|����r~�����c�wa�� )��J4LG.MC����Uj���A�!2ǥ�lqA�\��Zi;��;�1��|&~�k������0k#�cj2@l�5:�fWm����=/��ܰ�|�I�t=mpq%Ct9��<�۲188Ʈ_�h��k6^+� Y���Rju�cr��JP��D���<膕}y��%;��v��*2G��{�eI\�q��v���|<��S�0�(���V�|���߯����'��fS�Z���N���ɤ�Q� �sV�W������Gɉu��d�Ա�J�t�Z1�����뢁��&�*� �s�����g�(�T��Y��<�'���ktnǜZ@Nsm�?j���������b<P��ӊ���ɬV�B�ᰞ;�j!	G��VF�q.����\A� [�9d�hi<%�
p����ܙހ�����G���Km		�2S�Y�@�MO�PW&3KGg��_cؼ-kn3J�;v����ŭ�Ȯ��(z�R
-q�t���b�����L�vJ(�HHL;���FĖ��}Ǐ�w?t�r��"x`t�?݉4��xѝ��l��7�5a3�j�����ڽ�)I]t|;�jRh��PAi
f��ueppL>���ATx�k_sۺ/:|�mI���B��acd	�=bO=�t�÷���,���)�R�d��'lseK����׳Fbi�������g9Ɏq>���N}7�I��e���j�:{���~&���L���xQa���R)R�L�W�ں��@�+���yo��P���u��Yq{~F|G�$ϐ��)&�׈=W)��s����?
�hG��/��͍>}L��}�>�������<��4e��k�g�mҷ{�z/��l��Q��^
.`�|O�y���́���-�Bb{�z�;���zd�m՜�G�Z'�q)iW|�Ϳx����ڃ
��>o�n��n��!���1��:�����KFq��'�]�5�)�Y����H����S�ol��M9��;N�E�
�<E"
���%=FmH��T�5d[NW��n����fYė��pjݦ�5b�s�����5;r�ht��9�/�K�&�aW�٦H)�b�R��v E�%�R��pQ�$9�
��R͍ cb�n���>j���~�#�������cs0�����ϧ��W��#(ʵ+�+z81��+���g���wM?�He=�[� S��ʕ+}���꺎w��yϻ&��sF2fG����)w��fe��^�����"�㡔��N5�N�F� ��C�1"���F%���D��k"S�C!u���ڨ�v?ÛAan��H��G���|�{���Q��	�c�(�Y�J��̯��o8�=aox�p�*�Ht�u�FZ�_�7�T��_���_-=5Kx>D�0�A #�K~�7�����ڶ|�|�K_���a�7��[�P���ƣ����a��i*Y�n׮/9�	����.b�UT)T��(��<g���X���#G�M������w�{���?���5w�4��\�|=��MoV�@IYn8:�7yf�(s�DF���,�!�ܳ<��,g���=�W�H����N#C`*ɲ��ެ�	�u0Q(r�� �Y6�&]锑խ���:��4�`��(r=⳹!'RW&�X�\'����hM�P,p.�\U
lR�]	�T-����Sy�������8���Ġ�5��	�E�-�C�ehf ��^Դ�j �(WV�l��<`������	����t;�v��F;4w��l��EM�Z�`l���ۜ��k'Jg�j�u��Y��! �׃s^X��M�Pe�w��Z=���(\�׿�{����Z��-��֎(�@�aҖ{TۻwZ�^M��ť� �Ԅe��/�:��.rN7Q�rc[�b��]uч<́C�!��O��}�S��XV^�D�I���,'�	�e��5�� ��畹��>bS�*D[3��Ud���#�';��bU�(��&̝
&Ci�����{;���~�M��s����^���"��{ٯ|G�ԡ$��嘼�����o�	.q�����������G����_A���T�
KT��e�P,6T^��*�dj��n9 ȑ<v0�� v>�>��?�NQ�8.���VvB�c,>)�>���_����E/��b��Q9I�
�C#�ﲕ-�<�6�<hoz�!���^�n���M����;��sO���e��ϼ���?n��l�q��x-������
o�ȚlI��c���߲+��F�;VR	8GK���E,N"����.��;X�띦F��`z@W��̜l$�����٩^�	$�|�z�~VF�s���1yݣ�����PѾ����Di��F����jn%����rc-�u����56C���.2���?�n(!�Pu�$�̍�
�õe'&v��w������}h�� �/�{�W��gϜцPQ▒��J����O��'b�<��P�����G���FS�G2�l��X�Dj�u9��h �G����ܖ�x�})W&:��I�?7��={J7�.�S���x�O�Μ9�g��D���	�́ڐt�p���BG�  Y�SM<����u�v�}Ö��l> e���cp�|N�{������݁D�G"DEzI&�\J]�=E���<��~���|�mo{��}��*S`��hȢ�V	����5ᇰ�	��k�a�����)x���|V
���>�����'��������.�N����)[\� �<�s^w���8g�~OgɄ��]Y�0�������p=J�[-7>�	_����-��zT=<���X	N�G��6��v��Y7ĳ6�kZ`q�޽�'�2�pg������40�{R�2s�,���zvn.5m?`�~�H��%��q�Vdxd�� �o���o%��eu��'u��zGD/G���i�I%I}H&�#+���ª4܍�gZ@c%�=�頵�Db5J��
_����<���=�z)Eƒ�8_CV���^쌔(�QRN��8������/����g��t����s����k��,�.�*?���$�Ր�*��T��и��������&  ��IDAT˵��熍�	V*612h{�F4�z�h<8�iX���́ ���UeB�6�_��[�m����!�ƀ *�!ӔŚ)�����e���!{��W��Hݮn-J�R>�����@�_���_y�+|:�/FsEi�H5Y�ndf�An�@�n��t�Ĝ�xKMK[ҭ�A�~��O����}����=e�
�� ����yAU��m�ϫ!���}㩧�=��<vO�n�F7��[}�x�C���/��˻��/9v��b����( �$�|���rS��Pژ������9o�\]���y������E�����7�x�F+5EA0ȴ2|�y��9�; '���R����kK�`	������WW�Sy^�P-�X8AW��J{67���`5��9�hZ��_~ƾ��'����;EI⚗|ORz朰Y9�Yc��v�Q]ęck!3X ��}���z�� 5��C��~�M�����a�{���r�/���E�ק�؄���ۏ�ZlYc~�F�yC_�x���v,լ�)i��$\_��n������,�E����8��:;m��8��6OQ��M-��c��k �LL���!����m�����#����U��Ԝ��?�ȰQ�9�����=|�-n��v�gm�=�����T��!n s׃��-�	��܌�&�#��E���n��M\�0� ���=�r�?k�y�{������n�M{�7\l���=��3}�u�:P"��J~.���ؑ����*��R��VD7C�wq��xRM�պi!�B�9J���?C5s��K� չ�!
`%�XN�d��t4�rT[L �k��0�������"���9]f1e��#mS���pD�o�Q� �<A��y��ne`�V�� {I�$NQyX lr�����0 S�B�ҟv��"�'���#����w�����G_e1�"���xm��v.�(���4!�R퉳R��Z'ƺ�vPF+�j���I��W���.Xŝ��y�9��._�鑩Ȧ����d��62J��A�.-7֗�-��Ɩ���m�t#�P�g�#�_C�r����2��e��&@��GC�;�ks������Ɉ�����b�0���FVA�h��H.�؍,+"�����4�b��Ҷ�Ȣ�Td��;�#x����ԹxӴ�B�>�nћ_� �B�&*1���I��4M�w�i0B�Kv � /SQ��n�iJ�����f�. y�;� �T�8W?�z=��k��&�w�S�C8���Og�{8N]Ft`��e����(��!��gC�zii^��v=invU��H���O{�_C=�J4�l�Eq{�#�l�^��ʢ1p}��=F���%$�_`6Tp�=����G=��'˧y����<JRhq���JC�3?���G������\'U���GJ�|ߑC�v{yyQd�A�ۘ�UJ��l��jh�u<����;ͷ��l�KQ�ϕ������_��c��G4�����D� xR翯�̙#`jvB��S�̮8���%sSQ!�a��u-MTҼ���۩���#� �jO	b��Θy���.66|Ұ�� �� �.�w�����^l//X��,��;�eOp�؋�9�,���	H�r���_E� P�	�pN���Pј/H����*{��w�o�_! _����ĵ������'Hz���p�yE��%�)Z�#�`�������p"��܎9b���UI��TJ�h��K�VWs�0��wL��e���nů����2��h}��.�����7��~����6
��(�r?z�����o�����C�����)�r|2�fmi��+6L���9�vc`G6�jطn? ί�UID�6�ߣ�<�S�-+�쥱|�~�/G	�,i��t}Kiu��"�-e�W>v2)AZ�E�\�.pNn������^~舭/\�n���G�Xt!����	@�f�w�4���lQ14�T�#���jY���:� G�{�O�~�?�g>���E�4�������O����Q�hi|��(3��q|Ŕ�S9����AI����PqN�M%X� ��������e�W\st#���0�<�d���Х����2O=�tp�x���Y@ �QO���L��F-U5>*Jn��5s�)��݃)�&̄�<�TC�:Gʙ4M�ȿ)!�-��w���2�BF���S�=��F������V�$��q�9��1�ZwE�P|���=�7�~�$1t͍~�c��R9e.~.���L�m�v�I.9i�u�E9�^qPZn�q���ƅk�=�8`���Gm����ٴf�������Շk�#�4�Q�;�V����Qm1��*���d8�I#��ah��N�YPgAц�@�w��d���e� ��:�������^��V�5��Nk�/R�miVCc/s�b<_A�ӞdE
2Zp)?ΆTZ�^�	3hѨ-��v��Ev!���t�����:MZ��{�������b���^�\W9��ȝ^�k���j�j>�nPfz-���R� .���h e�d��%wr��dr%�M�mSf�N����9i��ʶw�Lԩ�ȚW6�� ����k�&M;q}�^_Ӕ�Y�H��Wp�R�+�8���g�w��ū����H ʞs|p �����˶�<Ϭ<]ȋilWQN��5>��))Nq�u�D�)7(%M�B_XY_I�|�68��˺��O~�~�a�� _0BSW��c��ɸ3���'�$�BWB��9�sH��72;�ri3O�ɒH��<�2ѣL^HM��{����~�W������f���ٮ]Sҩ�V�������[:��N'�Њ��Yy�����s�DU�&L����b���.�v��*0P���!�]�þ���b-"�2�6���XN\�z`�45�F���@�6\} �[���3�^eޜM�6>����������X��)4$�uHA�6P�>�;2z��c����"�z`��R�O[�Ü{����{arCv�
ϝ`��>'m�AK���/��\�O�ď� _��]�%�J4_b���W�C�c���^tB���权E��Fe��س�f�.ؙ�'�ֻ��i��>��W%<�A6��Ɠ�~>WN�W&p�\��n?�._����2�?v�,l�V+�x[6��j�����4����-Ŭ�B̃��I���C�&�,1�u#B�B|�Ӑ�`�׿q	C��,<�ep� &?�=�%��O���w�n�{���e�����1!a^�^�;��`C��t�6�t	c�P��4>��,×�x4Xpl4D��w~Ge�,<
����w��4X��J�~���3�7wlJ�>���+�?��(Ι�|��f']��9��M%��{fl��F����Zp���9ɦ��S��{b#��,�3S&�A�"xC}	��R���$ҽ�Re�e�k)-�e�ؠp�s~��(��QfPw�G�q81r���_ �5P��G��pX�yI"�\�d�{A:�ſ����s�����&��H�$�����x��(���TԍA�]ٹ�)�u�V��IOpS�p�mݼɍS�F�Ǭ���T������'wٛ}�>��/��ܬ�_���Z� �6yd�u*ukq/�Z��SO���9PUF���Y;w�-8��`��%[!��Fck����51l�a40�"Glӏ�+e�GR���sʌ�b�������̞50˥h��M( DD�1�9{��;�`�9q�4k>	�y��8���|73mr�	��;_���m�Jv�h��#�ú��t{7��́S�����罾��ZLݲIp>ʖmi[.\��`+_O9MhY[^K:pa?(�����BcnPee���/��Gܷ���ն��&�)G�B�jS��������`��!���v��~�%߻k���iK+
Ħ�L��j%t� ��x�Y���ذ��TJ��;g�f��9�,�@��t �t�Z�l�b%��a�7�� #z����?�3?mo��7������	4�9YD 0�TP��&��>#�|��@�ms��RHӞx�]U#F\�lyq���.l�M���7��~������U�4d͝<y����2�*lDt�w4�ߝzN��I���tfY+$�����y}iJB�~�y���=��	{��gdS9���I�����$5U8÷��HY
^�5:��eK�Q9h#�ɺ� ����	i-�k�߰Ǐ�rTv��3�����9�Қ$������$ �e�J��Ay:Ou�H��} �4q�1�?R[��>W���d�T�m<ǟ��_���ɟ��{MLnJ�H�TNɖvZ�a���3��^/Ue{]%�۩��jQEɅX�ؼ��M;u�N��ޗ�a����;a]��6x�$�Ԍp�҉���&��=�Z��g6v`��n�����B�O%쿠����c1p� ��4K����^x���F;Z�1"#mG�~���67���t�M���ݖ�VDl�����I+
}�6o*k�i��#��͓�9e�^Ss�٘w��$�8:=a���5��_�|�v�c������V�a����$�������B�l����Gɛ���JQ;��j{'���?�1��_�����C"�S @T����ӆ�#*�O�|����!�$�x�,xʾ�3?�` �I=K��(t�)��309%@ȂlZ��@�~$���ֺ��\u`��#��s��\����<���q��E~@�_#��&{ʹ��8� !#����C��(<��R�x��Ū�\�)��o�uљxˑC2����S� ����s�Sɦ��?�0����h�&7^�3�Ó�f�м��7���ߔ�!�g~�'>�i7v��w�K�B����	�Db��U-'��zI�����ɍ|Ps�i�Jɾ^�N�{wЍ<�7��?�
�z�%���7��z�U���I��MXmj��RB��]����ىS��`���t���G��_P&�2/Uh�j؜ȣ8�>�v�+`��-���W��\���&�I�KE�������z`z;x�"�km���9X�M&R �����e�K�U� �I��|��vӖ��y��2� �A�WS"zQ:����3��.�y~����������3N>O�p���(�Ȓ~,����4�Z5>��A�@�Es���/�����z��g����Mei15� ��[�~����ىW��ue�X�[n�+�>�n�Ѫ�������+�����=����Wm����U����z@5/���j
j)ڸJ�Jd�,l:ޯ�u#-l_V�#�r��E�H.P�m�
illA�mhxP���Bj�g~��׾�5�\��s��9��<���d-��0���h�!��. V��(�'��Bd2�$�T0��1��+Y���@�8f�w�@��P����<�D3�ɧ���F����-�I�@	��e�~�T�(��z��+ޟ˻���?p�s@��3HW���EЍ�@���>��Cp�wzFB�T���
�Q1����c��?�wnԣD*%Ͷ��)�/XgdF�3��W����</��޿��_�]u[M N�=rT�X��܆���x��K
���-���>�����=�ÿij f�8M�4��/�"{-�E��O��.��91~lhxD��z�rcǹ�B4<�qg���mW������E���i_��)Дt�చv˕hP	N����D�IՄ�vz$�,'�3�3�%���t���������xݚk�썯�_���3lc�O��ꂍ�'n����]���9)�*x��l|z�-4;�w��RM$*;�����^p*��&�����DP���"�̓��:��ʯN*I��#�2�B?�r�$�.*���c�ϧ�����n�,9V�W�z>�]Ċ;��ɾ�Տ�0zE��x4B*X���rJ=��e.]]U�i�I��zù�)���*3o�ccNy���?`�����ͪ�ݝ06:��S4���19����Jd�I)�X� 2����LN�?r���۝>��Lݚ,&��1h���ǚ�h)�R�9�w!bc��H�� s~p2"b,Ƞ �T6��`�~u���SY�sR������ ���ND��������,����"���J����}�=�\dz�*��� ���NX2o�O��<K�����D�Y�  ��;9��P ��9�WeC	��h��t�vR��{�k_�����~���g�yZ�lj�Y'k;����̴�1IF��2���IBR�$G���<Ң+�`.�_���9{�w�ʝ�{��/8H���;����HV�H�A��|�]u�v�]9�ʾn��uƇ�;���H �^m�1f��kt�jl������e�,�!�k$֠����s��=N��r1�I7lhx���no�ܪ�brH�����3p�1=	�	���S��\�He�cJJp�}Y�
��@�AF�{S�R4��xD'�ίM�ڊu��b	 A�(5��R�0�����i�]�(����AհB��T��,�l�T���t�rXW�c���;�J��(�Ԏl���=�?#c�kf��Pd �wBT|ܣ�%�HV<�v�dI6� "&_|�3_��|�v���M��#���);�V����T�*�����Èǋ����o�馦Gf�+hڐ��ޓ�*!0�νVG>�7�m�п�_�����G5;\����-qoQ�XY�������A�^ʼ�����ry�s"��� QPp��b�T��ڐ+:��h��?��O����na���e\]h,~�P~40 �>H,5������V���X�,֌h2d��.sw�����ֱ8�<�~:�u0����s���9�m	_�)��"�;FU���4;R�'v�o��s��?8���9���g� F;Q�Z,��o��,�QB��C�'��)_�;r���<��G�k&������<�" �{"af^�7��_��$��V�¿�W�O��?�@��?G�/47ĳ�SR�x�u"��G�ްw�]$�Ȼ�)�P���@�̞)UUV�g}w���?ng[s ��aRҨ�}ǎ*�z��E��]8��t�q�F������1/�J�B��67�.�n۩r��U���?D�v��݃>��EY˪Z�߷�����5{��K��x�$2-$�(2���N:?�H̙�Yz�D�w?n�ޘ���u��F� z�3
�jϤM����Z�č,��$	�7��_Rd��6#ir������D_B=͕${�{��د��/��ds�\�zD��񇌢�MEJ.���ϵX�Ndu�C�4z.�nk�mg!bSS��i;�=h�Wd�@��W��`8�\*}�w����_����g�������h��PM�����ۯ�;�(O,8�\�����D�l�z=J��s�Ĕ�ڌt��2�����Q�^�KS"�	����)����d���eC���{xN�!��g)!%�L�Vϼϯ��T��f�W����SYYm*�@6��'�7��������7Ms!R�MI��Զ���!�[�v�+9�NS,�B��Ȗ�!�������r����z������;:q��ƒlbG㛺1ӏ��hhr*Ȭԋ�l�tl�k���f1o�<b���}���ۉ3����c��Ǜ*�����V[Qs/I:��[��*���hQ��9���D����:W�pc#̓���:5�(�X��,��m~^�8�^~��>*����J1u����6�,_���+��1�6垒xy`�N���t��R�~��L����/��h��3%�4��1ǰ����d�r ���4�{�n2��\��N��H���Wz}��z�R_!!�����i��7��Շ'��@����ܢ]��>�����KWl�m��ރ��*�r�O��2bM�[~�Z��(Ee$���?��æ��|G)	]�f�b!��CZ���Q��8wR85�#���?�G�Ⱦ������Uqx�|���d�%Z�Q��~���zT�H����=��RLB�7�_y�� d�Fō�*P�#��}��_�yQR%�S�r>/�F@I��(���_7�i4>�3y&2իL!PU���b|J~��0�|n���="���Y��ڰ�7�$�R�Q�cjT/��+X�{���hW7ݯ�g��@��U��Q���=��C.����>����{eϋI3qoҌ�zu��F�n�)�Ͼ��C D	?8��
�	H�?\����G,�:�#]r8�Q�Z�$��;Y
0
�_	�8�5��L����0ɡAi^ט��4���כD	����7����?�/�H��MI�b/���I�_d�wT[{�[���b��tdT�g��z��=��/>y┝>��������۵O�zs��縵���������e��A�ڵ9���A݄͢�6 �^ut�w�mV�[����:}�E~yPS����C�b{�E9���x�^���r�J����K����yn��)��gibR�q�\HƦ��
esbcݵ;z�v��ö2Ն}�P��A��b����s،�}8���������dI�)p�.eC����[�o��UTQ*Ţ�t��@��'!g:���H��a��I�R����^����j��<$c '��l6���*Ľec��#���Y�M"���~$���F�0l$k0`�+sA!�R��s��'<8��	��d��ج%6ߣ͔x��R�;���V�x"��7�pVٴ�ł��LQt3qJ�`D4��@�|��9����?';���D^�9�焈4w�i���ۜ�U�m3��D���!���*ݝ$D�e ��\�!?�'O���U�w���u�����ʯ�]n9�ƺ �Y'u�V�^^7M-"����eS{g����ęS������I�tG��\Bc#Zd $�|��Ρ{��c�A%�N7�
�2:�{�:�4������M�%^�_|B�5>b��^_Sö��&PX�E��)y@kK�h7���<-�<��E�kI9	,��ċ���1�<� |��������9��Xh0�ii�q��i�l���DĻ& А^e)�I����m	 `*'��ۤ+ٍr�Tu�,u] �����i���$�?K�O20%G�]߷��?��ib��_�.+�[���S���`�&�=%q�Z*��1�����};E�Y�t���i+DV�� ����c�W����s���}ay�^:u�.��ٞ���A���T��h�A	�f/���Ue��;�E=ˣen�혜��n��E���g�i:im�ɥ��wf��6^���k���{���;w���Mё��������74FI����)9D% �Vf�_�}� z���!cS��[�;��8>�	��?��?Ӕ�˩Z!A�����:�[Z�yny~���_������ pѤ�Vt�汌�#fO�8�V���Z~�����{��)�'��� ���s�1����l�_�ҭ�q���ůT�&�O|����At9��4��^�>�XJ���v��f+KGҟ{�I�F�߿{ϵfP������;nW3
����Y�|�MO��s$�ɗ��
͕</�E��/� �F�R^�wc�3x� ��H��H�����C�ܻ�ͻ�Fۊ��k�� �#�M���|B�D�*(�v�\m*�B�F��L�/���x��>~��[�n��g�]l9�^���r�qсc��©n��lw��Ξ9c{���I��ڢ��\H6%�/��</��7�]q����n/Ҧܸ���ͫQ�^�|�b�����I��g�31A�!�݋{1��h�o/:��1�N7��ִ7�@�e������{����Ң-\�d�z�8�OGzV�&I��f8������r���]H�I�"�Ѷ�(�{f��i�����k��d�=v���`c���q!«�tzm�wO�<c@`8we.�:�l���j����$@���4������yM����f���\dfXy]����t,A�kW����[�qC `H�y��uЁ��O��>Y���!�&�X���"�&b�o,��8�)B$a�X�S3OM|Cľ''��T�H�\ۨ_cҺ'\�����р���������~���i��qĨ��=�,���Q.�ӣ��$r:��F����i���`��-��S�%-i�� EK�܏����_���?�1��_�%ik����A�7/A�YZ����9kc�RȰG�Պ�qv[�H�T��H�6�N����ɓ��º;	c���{�eC�<d���KV`F9��1�%��km͍&���&I0�[v'M#Ⱥ��;��^�C�^_���y��5��3�O���_sws 8|��EɢՃ��x�A9� +]�P�wnܚ�%�x����F����Lؤ$8�͋���)ö�+���F�q�tg<��@ɢ��fM�*��5'�u�,��d'd�751���*�/z���ԖVB�LF��N���v:��Y��m
eFg�na�UP@�����Ȯw4w��}���@}$@���2,E��U��*��Ht��H�BA��G�1v[���OI���yݟ������:}��(P���v��;�������k��H�	 ;,h�1 vЏr�:�-�9	N�,��$�~�HCe�K4����lcȶ2y�M�.�5�_�����M��A~�<�뿲x��ꪬm�� 1hI��C3L�:�6p����C���(���5�Y*D������9:�3�=Ѣv�<����߶|�O��_����}��r�R`�@z�~QH�E𾰥��K�2ek��}r��r���>�_��L��dA���ܥ��!kI��uCu����I��?w� ύl��a"_S��<��{�IN_�=���>}V�[���Q�{��s���ٳ!�OeǏ;1�XL�RÐ��M�缵���#ׂ�VwK���1��l1��4�1rrqA�U(�}��=K��^Ag�%f>�rsb.�3,�sC�}�Ԥt+�<#�C's���)z�1��zPs��/ds���˩dN֗�j<�����]�����~��������W�l</M]���<��ғ�J�N@'!�N�ں�?4���㞃���v�꜕�6���=b��~�^�]��ے��wh�V}�ԫv�;�����#�����k����q_/��y��:�IGzJ�-#����?�ao����Μ:�lI�j�UF�!V������N�t�1���TN+���R&r��Rs܍nPo���9f����p�8�J���v���er��{�w�-��vu=:�r+�Ľw���e5��V���b�'	����5�������$sOH�������X�wJR!�$�HφP�Q�F��~9�cql�ێߦ��u��fg�JN�j���\K�V3�n�5�4�4��y�3��5R�Ш�č�9A�>�R6�7�wB��8�O�I��X즱i�;��.qeΞ;�L�s��$�<\��s���~� 9�f�r��EjlN?��Nuer� /F(�17[!�B����"��d=E-nz5�D"V����z1�ܻܙM�<�����9�W5���~C��	>����+��+�ͳ 2׳W	hIkbp)M (��K�l�4p��65��]�D�Z���A�j�\�=�~����X>]��r���d5@#e崿�B 7�@���F|�As�Hk�T�����%��Srݲ��y;;{ݞ��?h��`~�L.#�FPU�5:/�ڶ����J@��9�5i��)ɕ�%����S���r�I��j�l'..����Z��V���ÍȒ�$��� W�"��^��M	h��Ee�
X[*9���{u_�4(�5$P��Ά��d=��;H�TG��,!)�K�t�w���8^kj�3l}���x�8l��VG����ڝ��09�
On#����65S�W�R��b�f����5d[O�R�jB��߉{� K�����}�}�}ˬ%���z�Y���@!�
�?$�a+��-KF�-/!9Bf,,	�!3,a��0@h`����u���5�r������=�97of��?�7Օy﷜��<��<a�ƭfh0�/���Ͱ��c���vaxJ�"��f_7ش��y�'�5�tCF<�m�]{{�_��H�s1�ЩaO�W��ܨ�=O��F�)�Z� �T�iK��Ysz6W�m>~���G� �9_'*��t##5�m-��f;�pҀ�S�Bm}��2;�)�F��J���������`�/���d#����e?���<��g?+@��Ձ\)�|��]׆��Ø�ɂ��&����Q����h�qXI����l��'OT��X'�m"�M@AM�Qb�fp~>��P�@vOU9x%���_�̜���/�{�D:��ϊv� � �T�:?ۣ�?j!�5]Z^�}�~��e�q �?b�ҕ���V��\��Z��۪���;J��ص�(î�����/��].^K�>��x��L��CƉ�e�%���Ie�k�3�L�懔4����D�{w�����c�~��X.�]�>]��m�`�>�W���ջ�>c�24�&��fZi�F{����� �:MN6��|����o���C��6�Y�m��m���wX�K�!C��νDFn�&G����*�x=�����4��%���*�GJ�9u�/��wV�2*^xh7�i�����TÕqV/��(�!���f'Lؠ����p|ꐨp�F��ɞa�=e���R���d����I�!3P���|�� ���lF����憀[>�e� �LT�KI;8-x;S
���ӅG��V��~�$�[��$���$ѓ�ݚ"��k�}g���Au��#�,I�3����V==vX��S� h+�؛� UJѫ�	��X�DIy���:n4�����@,< 6E ��t�Q��;﻾mǹ�)���3HP~mE^.�����{� ���Q�'�0��O������S'5�4Ť��Bq��g����W#c ���-���:�y�u�Fy&��:�����~�C?�w������h�z��m���\R㧔@l,tY�bN��S�"隬��1�1������#�{?���k��߆�!ۏ�lc�TIF����6v٤X6�cS�$�))t��+�C�l�+W�:��` g8��̱c�nꈧ�W6���(~�߸B���Z���Gc�ѵL���V֌��Ē
�3��|�3}ǉhr)"y!]DCM��|E�<6G�BnL�j�6���N��U/�ies.+��#��x�N�PJ�s/,�r+��'� ��Ne����{Z�z<"Rݘ�t�y]�%�Pj��럷����=]�n,C��S]�7b%^�H�~ =��Swu�6���4t�pa�	i�^��C#*�V6%�ޜ:�i9��Q���q q�/�B!���W��ш�k>)z/=R!?WdN`�U~nN�����-��)g�l�Ϳ�W.��̦�E��
I�	�s�q#��i�d���L`,v��^3v�2�D�����N)'��nŦ�l^�nZ����b��'�o"��{��_���+��J�27�-�V�K}r{� �\��Q�KƝ��5�]̠\�q=�D��Iz��N�d ��ݻ�G8�c�FP�e���H�Ա#�d3GF�D/C��ڵ�h096*f
"��ޓf$�j�[k�O�p��٠F��b k��1<���i1��G�RW�I�<�,��Ԅ��m�Wu�>���8�RA3����� J� � ����ؖ�iD��Qf.�]c�c���;���d���-u�X^� "�os�FF�cj��y.�'0?x�^���/6Ä������{ [�����S���Ï����_Y\�:{[ w�ژ�R��u�N��v3-����l�J$�,�Uc��4u��?�S��sgg���[�����*��a)��X���8�5�n�n�d���Ŗ��|'k�xD��<Ks�#LU��4[w
�����?r�h�Գ<����I=������)z���p�h<���Lf�N+�����G6�j��ɲI=lo�&ё�p�xfF��E[���-U
R��tuݫt"#֥xػK=�E{�Hax�4!ô�
�e|j,��������������� L�&�R���;1e��[�g-�V3�����cy�3�3}=a&?���d�������������eS�oldT@�󳠖�����l؂�S����y*��"�)�79��M�*l�����XT33�2����s���Ģ�1. :�S�QR�[}DQ�M1�}�V���5��k��u���)�Ƌ�d�� y�&��E�'7��[{�Pc��L� v֞�q��eO����X�7p:޸G�X*��>���zx)S��_6.o|��/~�_���?��r��-��������$���S.r���D3��c=u��{�9(Jdמ;z8|�������� ��3F9m�����+�#��*�������FT�<�M"��l)@�B�r{K��u���pb���$�����t^�_)/�6T��W�/���x�w��f�+]���Y(�U�IN@x���4ً�b՛�ޚ���mV��f�����rk�V��X)¬S�d����,5��� #��؄vX���6XgH %v�买�Ȇ:����ͣ��2iҊ�  S�i�O�E���=k!y͙Z]o�f4h+*kI�Q�B5ie5stv�z�)E=�Z�ϻ��8��F.)g�-l�2���iʆ-s�N�5�:/9>��ZM�r943ΟLY�.�����:Q�F�lC�Iw��юB	�4��m;N�?_!��rN�Gש�����>���m�|%�,=�v����N�;u&|��WB5����
�O}�.�r� ![�.b�)�8�Z�p��iF��TO�L���ko\�Zz����{�.N3 d�������Urp�ܔ�'�K���m������� @t�VCg��vRDR|�����u���6"Rak@|��\tw?���O"�W�~�<4;Q	�O�5ߙp��e�>�vMv�L����*9y�t��*f��i,��sg�	a��C%E5?^�^ɹy~��'&�.rtt�>�(�MD �u�ȴ��k�oyʵ�<b�����r��0_�ݱg���%L�}��YD�0&��� �`��1�h����e`�F~�R��d�/6G �d��WQ�ey��ײ������������C�~g7��#9���7Ĳ��Ge*�Ҩ���E-S��46���j9�^�;n�?
k���Wq���Ӡ���6[0'mmeZ��ر}˞wceA����bخm	���.�~j�[�vPK�Au]��3�Ү�H�0R�f$��V�/C�72�~�1��y��98H$��u��Äԏ�x%L�$��X��]M�?@� �ytv[��"6�������Ix�â�&RdO\���-��:>0�D4�#jԈ؆S�(Zꄢ5y�	�0irيwVy�Gr���m!<e���!��/�4�w%���)EJz��cL�d�&�y'O���ʮ<�	5���9�>^$)���d Z�%�UH�q��9�h8 ����N�����Ȍ�ݻw��$�9���`$ax�������)P�h��jR� 6��|��`�I��0��^��ʙ�è��:��������a�#7��c���f+�(޽}[�`M!/ݺ����ߤ�Tb0�DY�M���1-i?��|ϭ��F�k�$������p�����'�)"2Amt��l��n6n�qAz��s����� ��NRo7n�in�t�i�d�>����җBX��&�$��W�����ԙ��Q��J�g�^T�"�Im����"]��P�ڪ6n�y��U}sE*:�Pb@�� �uԝ5ۑTP���=E� �%6�QE=���w��3)@�*����=�F\k�(ܼf6���mTv���N�>�"5��F8ȸ#}��^�o�֤ Z��"�Μ�N�궭�R5L���#�F��𸺞�=���&�/�s�R��������8��Nש�v�>�y!�(%*�d�ʕ�����N�؀pv��%뢥)s�~�Xc4I���]7O���t�2���L0���pҦ��P�U_È�\�_c����m�	�ȶ�m���[�bK*�6����EDq �z���as��E��6c�a�Λ��m����)��XcԞ�w�t$6o�� ��t�`{j�٪�aD�bپs�s声B.�2�����T�q�U�)��0�Ty����B �M�d���܅��W�����?i}1�xqa��7�~�ݨ$�vݝ@��di8�΃�eW��Ι�pJ_`R���,�j�O��kߥ6Vt2y�w�I��Қ����ݲg|x����EsO�:�$<k�'H�)�`�ʹ���鎭��=�o�ղ����bm��KZe�/΅Ç��^�=��,�*���C�Q�Q��;[�>�;wV�O��}��i���׿~M�u�p����
���d�e��#`����J�K���k����j�I)�	r��I�˞��<�N�L���T���"{ى�xe�9���!+������0Ls�yMTAc�x�� ���/��o�7��Cp4�A7�q�e��!�6t���g-�+1��}m-�>m���3g$�z�0��c�Ç.����5;=���A�����Ϝ9�n7\�������7����@Fͦ9��f�>���.�B��)�@Q,��%2�a��W�r�3���pJ7VT�g]�6���·�'��^��#o��(�����Fp�BW-�*�����&�:��O�>��y1,������p��M-�^4J�(�����#����~��6�� *	H���
ψ	�w�������K�76|��<�����U_���(e�="%p����1�6�6�����f�y[ ��')&?�C����� ��#������=���K*���ׯ�~]="��e��D�s�@��{����n�{`�0�D�u?Fbk*J+ l�i[u<��
�Ͷƣ#c�b��1�D�{؋V�t�-���?�էNr �%�#�>�9C
�uKJYW�7�k1��R��6���/�	ʽ��ӟ�t��\�o�`X]]�7�q629�Ì.]61"�ْ79�.�t���D$dc�90,'n���T���I����w~���;��%�5A7���vz��>R�oAM_�ݺRm���My�������G��8)٦��K�Q��͸�u�K�ˮ�}�:̬P���pr�k#��2d��#Po�����C�il (��Q"���S����>gm'�gw�h�n���{�C�4!�y3(O E��,i��m�<D�r���밉��v]F���^���ވu��N�@�A��E"��lK�?����;���us����������n�&;��O7FM�_�sO�O�)Ԧ���!��'ʟ&��5�|N	Ј�ڌ36'�v���ks���$��3D���e4k
���>��{�7���/�FB����!�"��.v"�;�[��W^xN�o��m��ťXz��h)������'u�{VENUp���Htg��}p�j���!��>=�r�ə�]�hS�Ol9Ғ��&� �/O�0���u紋�����{+֣ccЯf�r>�c�se����Q�o�sRsҖ+���ژ�?LM�Rf��O���'N�e��#�p�G�"7nK�L"bf���>��r��1ҳD���������X�VAv����J�Y(�Hqc9\��p��D���i=��:ˈ���'c���8c�G%ʬ�{�d��J�Fi?_ �I��k>�]C�g̗���e'�Kί(������O�������X/���5��"����M�݆�~)[r�z
u�U��y��4�*��<s�����'���px����o=����q�\2�Lfۏ:�n�X/)�nf���Y���}E|R,��D�������;�廧:�g.��W�B"�	������ƀQ�<�
�X5�9H�FcW�n�#�����𩃚�~�^�� 9,�Dz*J���fgg�������/��-��oٸ�L�TL RD��7�4�X@`y��K.篋�Z�Iu��&rΜ&�j���`T��C���0	�4g�"�����	i;o:�Ρ�S��846-O[,�,
 ����u������c�%z�3<1Ǝ뜶	y��U���\�P1NQʄ�������0{v��$E���8IK��K�K�3(	�S�ITc��Z^n�#ã;��M)�Q����~�^ĳvN��mᲱ�6��I׵+劺��l����wŕR_R�����hI������?��x��o2}ߣ�NE�Uw�wb2�� �Y��M�˦� mb�#�/�G�'�^��}׷~<ܹy+���°��5�Y�<,z�K��
�$��k�6���Vؠ#��T�d��ͶQ������ښ�Ś�ͤLA�R��/U����y��Q3]g�#ek����U	;kabx����H�0Q@7����	j3��ŧjt�HK'E�t 4Re�������
���:ܧ��.�|�Din`s�ͭas�c��*ŋfS�K4N��+Жގ�} ��S^�S�7�����u2"�I����.ڲv�=�m"%6G�B"EߵgM@������A��;��7�F�w@"i�5j�����i�]5�P5�Q���L5�T�����$Ӎ�0�����
ka���w~��������(JJ��G�ҏM�� �H1�]��q����ڞ�=�n_=��ǅ�%�o�>�Ar�r�Е]� +����e�ܡ'��u>{�l�c���{O��g�9uZ2'$����$��n,��÷X�+ӓj���=+�)����"$�J�2{�
�6B
�œ��;V e����Z����j��d�ğJ�a.�(jY��Q�-v���ȴw�����}6��C�,�)"�;T����wdtB�w�z��Ŋ�y>���ȑ���x�p^%Zd�8 �v�����C�9���>vw�P/��կ��3<��'���5�)��^�⍌l��!/"�Wk8mZ�����߀r�1�>G2i�%��)�3 Q�.��"���N[�{O}���g�GE�n���ݢ�l�?�'�
�r1�G��z'55�բ��r� ��yf4I���i����^�K�r:��m�U�=�Mcܮu��n޺M��O��Ζ9����/X^<�۶�FJUs�ʡ�m���7<���%j����o����>��8����|���K�0���g����d���6�46L3<sg��'Ja}��M�����/�L���j�%��kK���K�.9ֿno8|��9����/�Fx��wRV�1��^�4n��H��%���>�k$rUr��G����:����&�S��i�V5�B�d��`c� ו4=�� 0J�}u-v��nƐ$Y�n��b�%o��Dd�<�vG�h� ��|�3�:<I7m��zD�zq�\�Lw�6���K���J�߽sO����8�|����97�l���!W�kb�q?�x�wё�}A��{�u0�(�>z �<��:V]�k�KI��lR4�v:Tg�H�p���o�H���lT�q�V��y�����_��o.q��ה�������ķK��(����7�1#�*�g�q9Lڨ"��0�ܱ�됈H�^����g]�h����}=ܼ{_���ڳ���+�)V	����V�S�t�A/z�y���I��~(�~=��:�Q��g$����=P��%��Nl�0@���O��ś�f%j/�����a��f�6/�q�W+��Ӫ)��s���ha�#���]��L<��$W\��H��j���`#�G����J=u���ڃ���b�WH�'PϦ�9:�6� ,F{1��R�mP��1���ӿ3�����F��D`�	�x7T�1��ɶ���(u�ɹ��=�s��/ۘ�I��x:��"��;�X�j�
G��T'M�ŕ}ע�D�_��"�h�?wq.���@81>6���:mH�T�u_�O�CckӀW74l��!*��]=�n��T�����NM::�ye��1Z+u'j4ۮѝ��hи�A �����Q�e���u9Ʊ����e�O"2-Qz5g��ۚTMD�U(���"�(^���b
j&pq ���iA,`~��RXY���Ub�h�sS�N`���R���}�kpP�T��{ k�}|p����6�sb	 ��,r,-,�a2o���נ�ϻ�+�=�}ܼ�A<�G��@��.ސѾI֐�Hu*WK
D(��9e��P4)Dq�(.�K�&�'{5�9x?�P�ESV���4�:Q�[��e~P^��i(�ݠ�xF��h���^�>��L�̶�1���s���ԧ�o�_�KaqaQ�TE�~���z[Q�均�(.jT:ψ�)v�KD����{�a�g6��'m�|�k�����X6�CץCz7�{4������f��)���;׺��3���Hr�`W�j.uF^<��}�;Qj,!vf3�V������2F�@��N"��h�c�������Fy���W[7�ś�R7YWS�6Q��H<sZ��<�,d,5�8�_���~��~M/�N,6&���e�E@B/��KG�&7���FZ��2W$�%	u�=eV6C���	�'��]�ɘ�CV!m�%��=O����gue�<���c�"�z�qx~�O�7����e^�k���(<h�y�ʐLM��M���Be���R��T5)���~�P�xs��E]���[6Y�y�O;^}��0;sƟ!�)���'��w��[H-[0[�`�?j8k;�:��SB�{�*C���0�s]Q}|_�T\�rqF��Px�IU@J�ӥ�KQLu�W\AdUQ���1���5�KJ����b�Z�����.�N%*x�<P���{�tar���φ��gO�u���|9um��J�FE`z�:�Q�^Y�C���)���ۡ�(T/#Yi����JŲ��?�Jx������f���E��֜N�����q�zΝ����D!L��C����,�[��L^��j��zWl��<���t*�u�Q��Ӝ=m�nl����S�b�]-�x�9��G���F&l��Ӈs�:f^z�y.�ȅRN(��@8��vI�ȼl��J�+���B2K�(=�>�(u��gϋ���LH�m��z�r{n"�۫4�aA{��C_��܀]��%u��H�Է}OMM��ZX�Ep��Iy��LM/�#b�!S�\���JC���bUr���M��z��`9���;_���{v���Y�U�E��c�%촩���M �9Z�\��<�4��Q� �Iv!�$�4���Ù[�Y��ю��DԱ�#�����L�������K�ag{S�4G���:�3dx��n�rt�u�  b��؜�E���yN��#b]�7��s� _�=މ�
��^Ʊ�Q���v�N�8fgO�\�8jNCA���W����4y��:as�O�@Op��xB��n�=�xU�tT�kkK������3~��)b�ln������G
�LLy�6� �]�� ��-m)�̞9�g�f�8��o��_�����]�'��J
��ҝ�zOz�#�aE� �D�֛�%p�����cf���Ϊ�eyqI���A-e1���	�B�$ #s���쓳M��w_#�.=r��9������9M���>� �8��r��؜��|B�${{�����6��3�7c��b�G}xE��ގ�ܵ}�>��p��	�2 j{6�vjN���8]9����mW3��|F`Q�sh	Q�O}'�������}�ka��Jx��s�;_Z_��0O
�u�8#��΄m�J���^�Y\�$�<���m����QA�FM@uZ n�뎚���7�j?�ث�	�?�}(����Z�A���^��f�j���<$bhB�57lw�V$|�� m��4�-� ���~��D�%M�_���w���B�eR\���Z L:�F-�����Ӓ2���b� 46c2&>?>��]]��܋����^�QN�O4���JLmP��io����j艴L\ �ƚw�1�������^W�Kg��v��VKROLL��" �k��D�\Pw����W^��|��W�1��v��Ͱ�L!xY��c�\������Ј�@u2�q���G6��Z�DH�?��.���`��pm�UDxo(Eĺ�X��h�fgf��&p]T䊐�2D�[,�S�,~�]��%��}�N�i��ߤ��wS����l;��H��L���2��?��a|tD��B5u�V�D��rު��W�Eح9�R-�Ā ���+ʧ��ڎmK[p�AY��Hf��;�M[5;h%c���mk�����(���d��$1&ݸ�c<D��g]�cP��#`�)L.`/�6�`:����Кtr��\!��n�JɇQ��y{�D;Ȁfc�1-�Z��P�&�5� ]�hSt=��NU82v6樎4p:n����n��8�3g��c�w�5����Ijyl�O"��)Jiw�:��D`����i��3�͆��a"�C�S1Jߗ}�F�ga�`$�(� ��'BV%eO:���\��������w��I�Ld8�㵔� }mNk�M�ua����� ���0Q�{R"ڽ����^^4d>����՗^���1��ǡ�{~��[��S��8{��d�x��t7�6�Su�7ڕzQ�� m�?��v����� o ؟�����{����.�mo�dh�>O�������V�ъa�p��#6�i��N�Sѡd2�$J���������.+K5�`ޜ]s��v�g/��F)�b���s��x��wvv��3+XSk��'��LM������t�P�ݿw+�8~*|���g>���7�]�]���ڣ �p<�UiA-��x&��Q'��26��30���BY�u�N��߻">wG�46)oj�!LgϢ�}��by���^�36���eC����vxy�l0Y�S�O��h+Q��f}cݹ���������nu@GI?�x���t�P�!�R1���Qpq�8
����֝ۚSr��KdȮD�����쨣Tk�s�~��FS{)��[��c6|<g���˗��矄[rx��nN��?�BϘ�5ӱ�(ځM���d�r�;T
������v�*�f��u�k�O3q�TG��Oo�i\��^���B٠Z�x�B8g����b1 ��s/hb���F�:�v�b��Y�Eԛ%�Nj�ZA>�m�T�^����/�;��F�G������}҇uE�N��2�Fo/��h$c�7#P "W��eI�� ��@�&8�h�AI�&]j��y.j�HQ~��E
pCK �"� ��K���x8~�ꁜ �h�/9���D��$'��ft��Yͅ��~[�8��r�xiN�[[uy�4�p����u���Y�''G�PȭU��ɣu�q�q�?��^�;�v���E1�I�@��F��{��!m
,~���Pp}��ꄅ�����C�Q�į��S=Z�KL�#����5�,Q�*�$�HIS���H����e�@�qp,0&�T���1}�p�m��˿�+����/O�Fp!E�����{a��cƟ9<4ℰ�ءݏQ�r��C�a}�&F'�'���_{��X1����:�	jv)P�ե���l\Vwͩ���.]�6��td�h��Z��(���q6V���w&�Y�]�?e�Ԇ�ݷ���${A$�,Ou��uyXT.:.�8�	�e�XC�PQ@��f
�����u�LtG*k�N��1nֶ�ZsG)ѧ��y�y���I���n#4�7��U=^�y�ω��X��5o���I=Ӥ�F����4d���>0Y���}�5�^T��O'��j&�%���CD5jS�����3�y�����@���6t�Ju'���Fԝ�(H<A��W���f!�Q��{�:"�n��gO��<v�7���J(e��sq>A\�kE�R��s֜^u}7[JIz�`tTz{M;��]�!PqU�bKM@G����@#����O������c'��]Xp�P����=2�'㰪����P�y�"�pT���51 iʒ�W���Q�&�*'��5��7�f6�iT�DM��f�KG��`z��(��3gf��I٣M(�ln���9�
��ݪ�!�C���%����(�����C@���K�ko�n߼�����w�W]:A
��o��]�O��$Z���zSs#��xG�t���q��moڎM@<7��o�w&���Gr����W�Y��o�zNǣ����=ҲD��{�-�N�@�8�o����Zkv^�k��w�k@b*K`OK2��26�9����kP'�V���Dv������i��?����տV7��)�󦱑r5֦�lu<��̪J�x͸X��f�/�x���8^�r%<�ʛ�������HgC'��������'<�%"���(ŞA�t�v�(��V�=;5 �u�S�7�|��Î<\�T/���^�c�ƌw�&��HU�e��%�|�T�:|,���n�E��0��D{� &-� �r�b���
bW�@����O����O���腥�=B�Ǐ+����`��8��>���tLG=dB����pd�x'���7�c,e��9sR��L<�_|�5����H�� ���c2H���G�uJƨ�EN��kݯi�R�'ΞK�Ќ#�[<п<~2�{�=��.]�d���������2FOx��yJ�<5-�|߻�5��l���zv?��Y���t2܇(s�n'Y�yv�y `����>�n<���BX[w�;	��pb�mQS����^���c��݆�xV�%`#�t�y�I6�1]�,���qx_�F��(�b�� Ud~��+�Uq�6��Y��(*�b���>>����w�w�x�
]��)f��Y�mhG��%`�\�
��uGBEgEu�7�W��v3<?w)\��[G^��Y��ˤ��N��yO�U�#�o�kazx���Np�9�~h+��1�XPT�cz~ R�tI��&��~�UD����E[;�Q�t��=28js�:�4�P�˩֯ec346�:"�Nl�w�ђ�g�S6a U�]��}Tz9F��V#Ķ�"1�m�'C��VV<�2Q�R���D(����V�۴L��ɨ�2E��
�kQ��>��2x������]�3��:�#z�����+�`�(�q۷�@@��BȔ5���ط�=\�+"�R�Y՗uD}*�,�Ӱ��J�L�4q�|d��%۴ �O3�hN'�C� m�dB �'��p��&�0�!��Tʯ�W�(r6��ޜ�Nl�]J_��"�4p�5����~�'e3�,�~�9�D)�AL��9m�Qvۀt]�[�z^U,ycב��=�](�p/�|�*.^</��c�e�H�6c�!�J�屍���:��] ���xw%���3!݊�|��^������n�mO_6J$���ܻ��fF�v��uϞ�^�JQh=�")��[��]\Z��vt]��;�䉓�Wh^Ħ"�
����_��ɾ��5���;o�D	*5@��s�Wh��]EK���f�M(��+�?M5�V[����n5���6�7TwHF�:Tl8��A��-����M�:O�C�i���	���5f�12[.���@�z�*�v곿�Kᕗ_��G���i������iA��"� ��QE��Ӱ��Jձ�:_.�;=�Ax�]���_���N��G�:��d�38����!E�}ι؅J��
�KC�?��#��F��dԞE��O7�<���:KFzQ'@�j��xv&���6�O���	�w5 �ؒ.�$���)��z��v_�ӋT=��5�<����B.	��o�����J��a�S;���٩�9)&&5 K"~vM�/xx$|��!Q.&?K5p�jY��
�/]���qyiA�y����8���z���kW����䚢ۢt���ϔT�@��<�IL����s6���.yn>Gx��o}U���,t�sP/a�3��_�#���pg9��*%�;�mƼZ��[\���`�ܩ�a�r���a�T/�@Gm<z�G��>���Y��m����QW\1�����6�^���,G��LjJ����p����޻�y�mB��U?2�� ��{�~���t��by' Iu�MO�|�D�	�$��7�	��?��a��\�W�N3�80��Kt#�k�6RI5&qpr�vl&"RDd���[�n���������_	���/��6��3|��]�C��j�ڤ�'Ð����+gJJu����F׀!\U�P��=��q]ן����oA�
Ĩ688A?4Y��dԭ	�uRoS*�wX7��Q��n�nLyd�,Pl��F���fcLu��]�P�^�	�&�������Jf�����A��=�/�F<A޶}�����!��x����*��5���9�N��샕��^7X���{r����� �&����n�E��u����_�n� ��G;s029�D^6F�~����e��sۏa�g��~�@���6ٯ�sg�{���K��w���N1�ܪDg�fS���O��/ ��-svU�Q)U=�v�ve3�?J���]���
��U!Q|�6�@��Ê��3��w�h}���&�} "�uȨ%F�l���̓�jH�`AD猷�ե��p��&�(P<�>v���j�����Ԍ��k��g=v�/
��nlb&C��j;��.���v�yb�ھ��u� ���e�}�a��e�4/�9��J�N� �hoڸ�㇏m{��I�o�%`GF���g_��l'O����;��ru)ܻ�M,���9��=wI��l.Z�N��"���P�4b��"�M�dc��fR�����/����h���U��u��8�$��\T�aJ�<{!)�۷�Hb<qv����	e������]��H,}j6�w���^���(.;�N�fFKJ�^�t�_�^�J�6m;Y|R��`�G���3�£'Km^��{��]�����Ԩ�����\d�P�2�QYQ�u_it6��/�$�Վ<oN=�jb��\�9�4QD���2N���k"��Pъ��W�\��m�f8sq6Tm�@�ۛۮL=U6R�^w�ukz���5�?�� ������?����B7c�`6*�T�CJ�&�`�&9��AX:1�O>�{�[7�Ȕ�Hނ��G=�K����=ܛ����I俹ƅ��� �6��i���0Tx�U1�oǦ���ĤhB]�A�p��	���e
q)��[�(F��b!:���!���i���z'�2D�+��WI�5����w�}'ܿ�I5��<�KJ!PҦ4 �fr�D-��oWN��ƶ�&�x�^�Q�j|((��Z�X��~jo��C����P�I*F�c;��k���*�:�)$Y�Dq�RRP��!��A��}R1t��NR�y�<+E����{���~����J��1��ہ��rWM��������i�ĪB�O�����r�p~ƌ��0���ݩ6p����?�س��P4��=V�X�Dk�ʎN\Ӕ��l��F�� j��WثK '�W�4�7uA���DI?�s5��t�˅�%V?�r�(V��"�E͠BR	9�
x�N6F �wtH/ع�zY��x�w�*�~��n��s��P�z�qa��M�l@�h�L������{�Ɠg�Nr�(f�hl�1�:�dCZ��7������~�O[uóN�טg�
�E��zTi�3�~R�c�X��;Ew�6}����ᓟ��t��
����GU�"5W���9�*�=jn���Uӛ� ��d�R	J��3�{iD8ۭ����_��_����>򑏄����j̔��d.(E��OlDż�{iϨ��鵜��)�@�b{�T��i��z7�ѣ�Ը ���t�UZ�\�=z�h����Q@rͰ���fw�s*Y�u�Fx�����/���&������������pb��j�	d��~�������~�ϝs��!�g����;�d~Ԙi��+�Q��E�T|��^y�u���^�j��H=���=�[P�.�v͆o��hH5��W�I�'ʼ�2�]u�R�M���n�8#*��L�o�/�6�[���k��QP �[�����ŀlu��}a�i�e�yjR5��?0L|��ۚ��*�e����7����g����~iaQJM������$$���r{1��%�݋��V��MC�fӏˇ�n�����N�
wn?��fȀ�(��r�����J���HF9FE��	��I���sZ��̙=�X�d�B�n��L�}��X����;����<��|���05R51��x�FOD�ym&;�R�����`�ZŔ��#� X���W?��կ�R�ۊ�#�Q���e3
�ۄ��ND��P�|L62�РP�h��J��w�)Mh��;�p�����*��ĸv�(��#	t�a(��Lđ	�ꫯiЙLT:l
��Q1I�O�� LH� ��9�#��2>D����gd�� �*ݟ�� �⽒ҥ�8��Sȍ�(��!)�(e��t6e���^z�9�{w�*����Od���h+bF�h^����Q)`��_������ ��5�E���!"|����;M�f�e�"��g��7�������v;�S�$�>���f�%�5&;Q�_��o��_{-�g�o(�N��#*���I��ԩ��kE)8?`d\+U��zil2�wdRuA��/<!,|��Ц��vN�����9^i���[�x�A<{�G��H�C6�K\.�(�0c�M#�v�b�������x��)ʎ�Ђ(��<	cCcatx,T
��CZ<�����ô � ��F�-0(�l�P�:�ڎ��P0'��Y�"�`m�c�:6jt@�;)�؜�}y3ȥ�wm�2��5�\�V��b:�c��`S\�r������"��Lxv��~����q����������}J�E�?�<x��o\��@�(s�l,!�ߡ���`3xs��JY�/�>��G¡q�A��H�-*_���m9�"���A\�\?z∺�E��QpҎ��3���E�7	�y"�Ֆ&�~���g��T�-�j�@J��ṳ��1=I4�r'��5���V` ��ҥ��9�H�]�z-���;RWHQo���Ԉ�c�=�qyeQ��ѣ�i\�����3>zڜ$�SJ��Z~��h�z��^�?P�UG��|1�uu��R���"
#ƫ�q�Rl�qu_�+kk�$&��aO���S�3����'D:�A	N��Q����?Q6����s%%����@��W��"��oovv*"�l��^2Qc�Mȸ�7U*^�N�U�L�,4]����؛`=h+��V��#��7u��T�d��4�u��ҴO�?�zL#T�{���ƍ�p:�vO{�0*Svm?gFA~�x!��_���/������< ������b��dR�s*����p''=��>~���|�F�>Y/͞�[���R)�=u=w���Hd��T���}��\�SGS���u�t���I�I�>R�P[�˳���	i!��݉F�#�ԯ����Ջ�C�6�Q{�'���=F`;R�b*��+@�0r'JoQ!7V��g�(���&�[o����/��|��٩��`�&�l�H�I d���^�<JD��J���#�l���	O3�1�Lpu��$,ŉ�������YM ���"�:!���"��w�y���H��D� ���uE�xv>�^9yp�������ͦ�y�1 ���0����P���r�>���+2i�#�r�7c����K��c����۷D"�X�:�3àc�YT��h�z��IR���;�ϔ��w��E�k��BK�% �x���� Y/�o�.(��g�����s�rP}>���4R��I<�M����<�S?�ӊ��a+�fN��6Pb0��a��[��
�����]��`�k�����Q\�-=	'O���J�0�[/�1�{D��6�zmW� #Ms��v^R���:�Y��5���K5*�ӔV���"�K[둶�
1ڄL�!�l��*
$	hB:n�M��K将cU*����|�l��*#&�C�)�^��l,>�	G��'�k�'�(R^�2��22j��K��єQ޳U ��=w��uύ��dɲ�&�����i�0g����<?uʽ��g~�7̤��]�`��)P��= ?��MO�Zw :��^?�	(:H�u۱�2�w��?k��m�{�O�]��6��Ȕ���y ��W=�U�{ꍺV$[g��h=*�%�������\_�5�!h�?g�Վ
�BL�u�>g���/���&"F���)y�}�HT��u�K��q�֬m���Qz��!��gΜ���yCg���q���T�9�����ZAvkuiY���+���톽ە���-���rz���ﭭM��?V<�
e(אY�N�hb�.�v��f.��P����z����.�f�����bl�*�I�D�ubs0{x��]����-����Uu?�@�X*l���֛7oH���+��G�|�A��I %MG���
^=����a⍍-�$7[��Y#��tyJX�1Qt��H���s;;Ȱ�F�xH��I�H,f��=�W�SS���А��p�^hʉ�\O��ֆxcm�2� �?�s?�Qr���X�k�3F��G��ݧ�.��
�彦���"L=�eN����̝:n߳�{u�F�����H�طc����(8O�7�zVZ�V�bte��������Fɽ�R�q���׍Nn��hE/y�l�� ���!;�=�s���M ��la�М������b
1�|9�kz���"�D�,@�ރ������\�lB���{C�	LNLk�3�8 l��(�wN��a���V|R�;�X8޵4�"�ɩ�p�&? ��ĥa�vH=��0D��Yuv�Y��7"��vp���u���م�*�4"���s���W����I�=�r�Իu��N���
A ��:��C�#���`<R���� @,��^��<)"����)�k�o�[�T��y�ׯ#��^{��p��y�+:7F���c�����(�I]'�f��הH
�
��8կB>;?��o'u�3�I�'�e����)�����d�a�\$J��wW9�P�i~$�V���|��C]����a�oK���_��_��ņ�q�;Kmu�"a^��S��3���~�[����Q� :%|�Sy-x�9���è�����O���~͌򉰰�u��ls�����9A��=��f��!���j�#�PåMF��Do�*�����s�-��lm�4ou)]!F{�@�N� ����5�g�Y9����JG�N	V�-�� �"Pܠ8��sk�Qی_�6�"����ý��c�I�Q&�ڡ�Ru[GCY�|uz/��~�OR���y�87%�E�g)He�����/���@v��{��{�b�h:JeF���(�c��ɫ���렛�9��!�q6��e���D��>Nڜ��a�o][�k�y7v�^9Z���.S��<:��cSeG����H�F*-H /!�HI��گ������\�y��%>N����ۧY��]d�^{H����U_>���C�C�a8N/uwǎ�p����{G��ҥ9C���ʢ��0?���-HJ#h� �Lʦ=z�P܎ QJ�^x�%u2߹uC�����*렙ftlB:���7���`�ٮ�w�~["��˳�������i�9�W�~�g��<f�n�샢�V��XD0s3ܼ~U{�?��������=��c�8Mt(����ٻᑡ������7�Nc-L���1�\������{��)u(��zө�G�tk6n�ˋ*ݹ4wA�= �x�[����c�p.���|�kwpzjbox�0��g��;{A�u���=n�,�*ѧ�xW(�#�멬�����U��Ĥs)R�>26�.��m�)*����g?���_��ÃF������[���wh�:��朊���\��qPd�삍�������f��B�]��L5�-9�rNܗ8�4���^�D8ۃG~cm�����º��>��ɳ�j4t�݅�On��}УMb�	��p�ê&mp^�|9��G-d��N�L�]�wx�ݰ/��)�ӒQAS��ќ3o�4���x��?���ƛo�^�qb���tZ��T��������&�
[#�!�_�M�H���`�e/�G8�*��+�4c�MN�ԷcW֦˫e�A WԶݿ�@��k2�����޽�RV�T䦢x(��t,d�!V	@qn"�׮]�3�]r�N6�SYSz��8 �^z�E�M�xR��&Wsq�&�}�v���ߓ&������/JR� �цs����d"QNΑơ�I�W u~_ۛq�Ð"O���f��(����bI�͸ln	`���x��ˡ�P�g��x�m�:�#D�_�#݌ ����:@�t��O�$�!M��xg��<q:,�¥�CP���,]a&x&�%K�O��^#�[[�7��R���6�j;�Pw�ej��'a����	I`�oRWt؀�xXzxKکRWj�\�b��I;'Փ�:���q0l܇�l�W6 g�%H��l��������M����t����D�@ ��v��oI���.�&lI=�]Oat�f����i��p�UW�e�7� �5�)�����p��^�)U���i:����gE��/�}*B�{�{���:��{ �(YUyt"�N��:��s��\;Iz�G��k`ŝ�������sDV�����Ĵx�K$�@�y�9R�,�ϒٌM"�%HNOj�; ������Q�J�}~��=��o���Pê������U��8��YP�b�'�M�0r̀O�����~ΐ@��76��H��&E��%IU@ߡ*2���E���j �����.�\�R8V4�Oj��T�	���#�<b� GU�q���p��Q�A��؞r����=也�ͧZ2��Q����ҒV�A��̻FIǫ�����o�Ɵ�,%Oo���J� �W�</�)�Qc�#*;���0c�Ƥ�S�(�k7���U�����BY͟|� ���x�{�aX�Y�;g����+� `|Ԁ0�����A�C$StL���S� ������)�r}<@�{���u`���w)�[�뤢y�����
�]�������m�t��#������0B.�z�~�RY�	u���l/����i/�x��hG� 9���KG��B� ��>e{�f�f��0�-�qUP7�lfI�ŞD�z|����RI=�"�N ��٠���M�)� K�
�9�k�+K@�"x�MRZ�� Bw�#,u��`Ti5�;�b��������yʈ��0�UB�~�Y'���zY��e��YԫJG��6�aJ�X��^���'���i8틺��6K�.�5�-���L��t)`��L�,Bd	�H�o|E1HI�0�\�NM	б��-@Ʉ�<���y[�Lh��y~uU�oμ3R���B��'��y'߮��M�|��Nټ��t�q=R�tR;�`W�.�g���\�!�(g4�y~OJ���|�������0���3��? 2�R��� 6|�	�2���,!W'���syǠo({��y
 ��ز�~�6ƔC`1��"V�L�C�w�Y�3?q\��O��/��g���ߗ��:Z+���&����ec��z����wc�&u�ݐ��T�nl�y
C����__�㯆n��G�ۮ���r�q�G����o)j��Mk;� qTsλE�G+Fκڜj�j�16u̮m��;�cc�u�E9y�̞��z�HQ�����܍FK5L��-����G�S����*i7#�+��ei�Ap;��I�u:uqG��6��=J2�������Ԡ!ˤ���+��&Ĵ̳�~��`�ş�Y��{?�u������O�K ����7&��w�^����.��"���6�_1��<���{Q�̀\��/�����>>.�=���]�鹒"�����*g�����z�f��!C�|;�����ܳG{̹��ѧ�[q���%q��T@S�����q&I5�ƣ�h� ��(OG���гGǆ�)R�ҥ����(<|t_Mx�Y����'TZC$��N9��ʌ{w�x��.�x����2 8�ݻ�N���υC�����|lw��<�����F�yi��2N��t�V�
��@�|Ā#Q�'�t�4�L�������!7޿F�?0�����]�n߽���̹�b5��n�������p��-E�p����:��)��:b����۩S�ʐ�:'yf���=����ڵk�����i��vm0Gbڞ��Q=s�[�Rb��D㎓>}aNvմVT>���yc��Xq�� k$���+�p]����h��c=�y|�!`@���fc��4������OVV��o�����忬�w}}ų�q�w����ó�D�.3K�͞(�p�$>^x��0�dj,̯/#_�/�KM+������Ϻ����S@�ۙ�{����k�����[ٽ�n�� ���#�.� ��l77i�����뚬��%�V`m��J�b;�;~^�xcJ.�] ��13�T?6Ѕ����?�:=@��ʺ��3�D��j�߹�F�����̒TN��\rj�a����(���4�z;��%�y�;z���xa$�(��$�ԡg9"ZL��sV��L$Ҿ����]&�<x��O�Q[ (u�L��.?�t���OJ�PG����I�(�_� E��ک��hx��˜��q �5n(ţRD/������Q�xS�p�@�O���y�`���@y&�,���qM�(�Q{��ԯC��r�z�& rJԐ1�ޮ�Ut\�-���4fP?蚛|���}�y�z�È`x��^	�G90..P�W�u��T��s�]	����"s��]���3��D, ����ڦ�}���mlD"���9m0�a͆m�怍�ý�Ր-UU�1lN�i͐�]hz���q��FO�M�Ƨ.ڨ�:�=6��z]Y
�n2�0d����b��&��q��3�I��<�9����
j*(S67�Pۘ'�u]N�hX��:<�-�X�fƆ�!�ݒKgsU4A�����>:�q
������͸��7�=e��h��>���wO�Of�I���gݖ;��28�s��N&6�ͯ�|��2k�&�꘽���d<��</(#������?A�R��~�>��]	��Ļ9T��Kk�,R{��Y�F�8c$!x�� w�� �������L���DvP�1=o�T�HEO%�]�&$עP�N!��Ƒ�9�alί�U[_���[_S�ZbNHTi"t~����6�����N���A��6+�j�?2G��F���8���o�3[��믘S�g��a�oܸ&��.j02&Z���u[s�P+ԕ���k��10��F�O`@%K6��.�K/�ܔ	���ƍ[�s�Ɍ3c�P��iz�@�KsƤx�1�{#lm��yy@��(��D��؃�"g����X��η��@���I��f#J��Հ� &�o\�h���t��3/}n��K5H"�`��i���E���"iq�P�ʣ$����;IɚD��Ȉ��ŸA�����U�Ͼ�T�|R��D:6�Y��kS�l.�<�C���k�|�4vN�<�G'\�p.<\z
ʺ^�B�f0��K��,���я���s����94�[����6�luT��I&�7�n,N�F&��^?�M�>�6g�kAe��{�R�4s2�<���"{��s��f"0�:�> �˄�zÇ؉��\2�"Ԉ����X3��奰�������Yx�Jc�ZGu$�ň�虓�U���o.���C-	��:Gk�\?�u��/ .u�9�P�Ji�G��I�K�.�B6|�'>�p�[o���.�S��� a���������Ec�X�D�RD���{����7<�yD� ���g�r�ҿ<7�z	p&nH���򃰼��o�9a�ىH������|��X̉Ɔhтv�߅�a�ɢ6i���<�g���Ӻ7�r}Hdq�<CM��XO�
���晉�V#�����	w��<|��W����8���q� ��3���S�kr򰺘yV6�'f��<"����DXT n��8(���P��x���GF��`�����s���!BO[�^f��8�dWNG�k�Օq�h=?VTz\:G�W�{]1pzxr4�?�_]3�-����3 UCd�Ͱ�i��&�|�m�����N)@75J����M7:=��Wf*���Ȯ+��E.
M�d�Nw���hZ&w��o���J��iA�1�	i5�D�q̹��kpk�D��eR|��'m@�H�=��{8ǧE�Cl�Wt#�g����4��x���ԥ�d��5|!9ϙx�o� 8�����u&�����.<#�x�z���컅��u�S����׊��9��}5��e㺹�,�c܀�����m�;8fH ���+�f��_}-��-��ٲ�,鶜gl�{��r�5H��yA!DB����,Ѭ�4Ao%�SZ�V�l$��h���q�p���}^SS��$߼}+|���( ��+.�I�q��H��9������xߡ��i�(^\�*Zl3��|lx<|�'?!`��/9<1\��n�zuE�b.��$��Ź�������̙�֛_�RZ���4cD5��I*��{���a�8��m�>�M@k�4�3۳%�R�KH'K�ŀͺ9f_���jn����ŗ^R*wv�\����e��ؑ�	՗�mliOKM��5k�ը���Wd��}d6��l�;�~�ow�A(��pUޱ�ܺ}C5�/��� ��ʚ�0쏏���pHOv�򠎺�;r�nԛR�{�6�:P�P*���ȹ�ao�
p���>Z�^�-.�J��}uqӂ"�tw��l|��'�;l1@ǝ�)g�"�	��J����ԧ¬�{�ձ�j�)��d7�@Tf�i�-���=��9/W��8f���£032N=�x�Pe���۔�-
���?fHR�b_Zt���6���qbT���cɳ�NJ&&ֻd0&S��zΛ8L�rk�m��a(�5�E�oV��5*�v�TL��n�%͘��e���|�ח�F�rb\��c?�c*�]]m����! C��t@����b���ggR'=OP{��z&j^���D��"�s/qL��7�2�����j &c �fVD�L�#�c(��R�)hc �ų��.�.�� b�]�UW5�,@�d��q7NN�ɯ�j0,�?H� �?�W�z[�Lf��,&>�G������&.A�	/�ߙw�I����%�����	��#e���3v� �^� {D-ק#�{��6��\]h��<CC�����4JbS�S5J!	Lf3}Z}v۽]�_�u�\���^��F>	c�55XQA�qbܘ�J���K#�0T��{_
�hLYo��(��,d�U�.XΙ�o�}˼h��P��[�w&Ǉ�ssgû7��fO}�Y�v��э%$Q��#�vCk�6�x��.�����h��0@�>J�u����9ohٞ�h?��U�lw��C/����Llj�G̟��:��$-b5����\��j��>D�u�m��1�F�m�QW���9MSasaWҢ9#y�ߺ��I�#ӇD7��n)�Ս�2�gE3��;A;If<�o����s<K��}9��������}�ϸ��%܋�]eR*:�?�~��(-����H���X���H�>�ak���y���C{�q��ͮ6m>�պ��9�<�t= �����YM�]�;��d?m-j��̆8�z� �����k�9`f�v��I���?��$/�0w�[}�T� qF���D��0X��8thZu{^o6�s��y9r�V��� �2V�ɶ�����u���Ӈ����< ��3gt�zdf@�G*7)u�y��7�/΅	��3�j�ˉ~ʥO{�`���T8q���Y��~����4�m�pl|H܈���!e0�D���sRc�լ�'8D�6:�@��ӵ�X�?鍧��}�=����QD��{������r7n^�]�n���	��!hg�[��);�#M=wlO!�KF�y%)��-ퟔQo
�7�H�,]��Qe͑�RJ��%�#>��� �H)��!��O�dW����	�ey�9����r
tp�6.�E�趐���9��y��:�ȏ������p]�*�����X�4��l\2(ՙ�����ߵw�Nٻ���a�9S0'� h�ޱxs�9��L���|��K��޳3���ƽ�_����E!zYN/R��w�)$��*��M�j����D��.�c�%�Q�(m#n#�$C���D��WaS���c=G3�����]{��x�����t(tL�k.��]��	�@��5��V�Q�A
�d8�d|"~���صhI/�ˁ�z62<���^��7�0��;�40 ���D%�������O�M4���6���o�& ��)
��P��?�cEˈvy'�a�a��8J0������I˹��.��5�&D�3X4ep�.\������p��U��|�5��d羏=��8M��g��{c��X�S��k�6��H ƓE�����)���4�����}�t����X��\R��s�^��VAz���(�w;�^����6W��PJ�����`��mY�ݼ'6#�%�˚:��t��l�m�(ʀ:��o��o���"�_��):�ҟ��ik��~6�E��]S�\2�p�o��S��33�+W��+�q�Po��ܮӳͱT��B��4]�@t$��Z_V�ƼP6#Ք��������G�wCm��F�)jz{\|"�@_=陶Ek"��3*Pz��VJ=��<Y\QDr��a{�#�H��j����N��v��J�t�BkӞ���U�����]!���X�G�=�RN�u�'��H�\����޳�� K�;鹻��b���vp0%��t��uk��p ���?8���K�r��^o�4{���Hq(d�#ac�k�Ш�4_�t�˗���ڛ�Jz_g~��[u������M�F���I5IQ�(Jr�3Nl�!H ;� �|
H2HHb3�V&�%Y6%J$E��Hvs�n.����ouk���=����M�c$H	�n�[�ֻ���<��<����*|�j3��	��1$���D�a<cZ�����^.��'A͠�N\�'��X�8"��7��b	22{�z�IS�;o�� 4h��IH�=ݬ��z���6@R���d�7���y�o�Mue8�5)�R�zAM�-1=@�N.{��y$%nM�T0���/���X�@���^CQ������T����Q"��B�4���9:�#��r������t2>1,����Kv��YQl"R]���=pHM/x�nK����L�`�t�&?�yG����Y�=ER/CY&�d�1��]�L6$g>���/�o7L����=��	YX��/i��l~i��� V�)�H���1Û���Y��j@*v�I��)b5l<�yrlR6�FK��u��lP5���"�J�3�����o _�g���u�Oa�Q��Mca��		�d���9�X��瞽��W*�چ���c<,�sxP�i��ɱA�����ϺoES�jj6�t.d���	
��J|�z����t����}A��K�l�$Fx
�:��/ �N!��~sy��H��Z���M��i`T�fV��iV ǖL�&R4��C"��}" (\$hoO�F9��G?�dШA�A�}�{.G�O�/yo*��`�T�"��piI�lD��Jg���F��2A���%:��XX,8���p���p�ӊd�,D��57����XxqV�U���,h��G�Ղ���f691�.6�gϞսໟ�yeOY�D�,Z�D��,���>*~'5Sf�@�r�� x����V�&�&��X/W��v��
 �d�-dF�67��{H&3��O�a#r�D�����`���ٮ�酒P�����9��0�|�g���L�b3ǌ��k/�B皸[�'�ן���q&��Z�ŉ���X8��kɄ̌2ϫz���8[�ah�>�C���@�����Ea�ĎNu�b�`����vn���_9�l����M���rH=��ɸ��%i�r�/�Z��%-I��7u#��P���̭��qr4���8���$��psvw���w&�i�m��-M���-��l!��v�D |Ӭ#Q~_s��к�9��>�f����@�t�f�V��y�ã��	R�ɻ]#�Z+2\��F����G�"Q�U�-�_3�:�Ƥ�W ����V�0r5:/J^]����L��7���Z�d�hn{��#��$mn�|]J�"cY�ttu�;�j4S��e��áC�v���M=�O�T|�+�d�]��X����̭���=���#��Y�f�QD'��oY\Z��;�����NP����҂�8Pi���H ���yrtR�d�H���|�}v�S���/ќe�`о(�r/�^8�ca[v��-ۅ]& ���x���&��x-1�*	������p�����q��u�p��*]jt�>88,�%]�>]nS�k�����
j���a\�0r��2�����Z���];w*qp��-vr��]J0\�v�Ξ;	|�0&c��5|����x��u�)/^���V�;�����&�	WBrft�&&ƂpTR^����~P��������T��)P�dl�&���`�! �j�-L��� *��s�y�AaDS�_|^UY�8������o~��ލ�Z_�Q���X#)����@{>�!	�Jw����}|wdm��6��)�uP+���f����Z_�xi��Kg>�T�zgE�ae�4Q�E�,۝ϭ/t0~�ՊK:��;�*$���lj|���:n0�0[�'ͥ";6"�|B�u�7�"4�AS+��a�� Ro���Oj΅Y��YC� �ߧ�H��g����D�e�n&�t7s"�{���{���5�0�}�ρ��`����P���适�,A����z�Cv��R[{�֐R>�ZJ�#���CB��3�,>΋s�o�g�����Y/����l�jF]MW�_�sLً�~Q�iwhfͻq��N�i�rͻ�쑁~��_�c���{��?���Ø(�U�R:&Jc$��{�)φe����v���N,}����ڄׯ�oF����������-.ڞ�������O��dz�"[׼ؚ:}�J����sZ�k�%��0�1� � �F�5^�phXp[�h��xh��e��~#�|�?֗�b �nrD��G�-ǯ��9x����R�5�����۷lϮ��5I@�۔�0�"�r@V�;�%��!�ȸ�h��UV��mz�����!����Y�6:`=���+��듩-$M� �Y���'�!v;G6����	�rÊ�ϊe���k%��z#̪�@я��h��r��;欌q�94���h� cܢ������a�\(���f���wY�z��ʾƧg�06d�}���w���gF�s���� �O��	喵�K쥭�xy~Ɗ~N=c�֙��mFsh���v�/wu�}�f�>b��6��MLF|�/�fn7~Ef�cb�v5���MJ���`��ݒyl�����C�*O�j��m%�D����f|Ӹ�]�{�~ Ƌ@u��g�|��ߵ��	��F��e�%|��(�9����UJ��Y�~�d�y�fqĖ�fXґRS'�Yo�`OD�r���ѱ��'Y~�"�t��+#��$_��Q8d�՘а>��t]�mQ��g��ȫ[;�I3�hݐ��&͗;̲���p��@�f�� ����}�<`�g$�UM�Zw��%��Vu�n�v�w�h4�aʺş�������: �OQ�p���/�)ftӤ�s�099&0399j>do��;q�%�����Λ�x��S�,���ܾ�L�Q��}�5���/l߇�?���jY*�r��ͅ��v����^�޾�
Y��T��?���OmqeQ���ߥKWe���pͨt:7�����c��u�� ذ�W=�M���_/.�	8���k[�_�����rE8���ϗj�7`����%I6:�Y��UI�D�:���Z;�]̕�Ӑ�= Hlu�!&��hUT�ziVq�CN{��j]����^������q�j��������e2L�i54~���38��e�w�R(߼m}C�s�&;�>���R��R���`�=�hT }1��.��5"�`؈��u�R,V?
��x'�`WP%���Zu�մ��<��UR�rj��	����9N�
�m���
������B9�,�f��E��ګ���W��y(d�S�^T7l����������x�q�+D�o��1GA���"TY����'��>�=0����Q�=�ܑ�a#1122�, ��s��	��#���@5��>_�d��6�p�N���?�����J �0����g�y$tLE�U "|>p����x_�t���g D|/-@�ȝ�'�`���?�βw����ؼp_:��9�,��ma�<�G$gd����DDF�z�Z$��Ȝ����*j]�"}���Ag��w/�٘k�_SG]ZK��&����Ϛ��c�ӕV��i/���!� ��~�����e? x�k�a�C�z(��4�\%6����g�����Z�F�Z(�"at�q}=.I_q= H7n�zE��r0ՔH�܃�~B���m�2b˗�e�8N:Ȧ����7����[��F�Do���i+:(X��U��p�������5ԕ܌�skU��|��ݑf�|���s/d<��W���q�G'���=QhZG�h��Γ�?F����j*p�#�Y��yDbStk�-��emڃO��^w�%+2����K���Z�ݨӌlٿ/�Oe�<@4��.0�"� ���ٖ}����+�+,&#ʹ0� +Y�Vs�ʚ$V4/�k5�dl.G�e��[�لݿs�<YS�E���<��������2��`�F:�B����6"gew���Ȧ�`0��x�mR���/�

Yj�����}�]�ڹKA;�~�<N~�m:<D�M:x�0���7�4S�y�I?�;v{���r��L�`���3gΪjB����ɐeV�1����-�^J���a���D�c㓲{8����}o��ZQ6?�H~&��f����+N�>����p�deD�����l1�T� Q$-�^�n��]�#G��<�|���7:<�{�'��/8w�L������u��U� P��|��\��s�����N�?]�����~ �:�����"��	��T$݆m��ڦ�+�d?_ΏM ��Y��輸o�̶v ņ�c���P���tʯƽ	qe�{�?��B�ˈ��/l޼5T&}A�����A��t�ܯJ)H>q��(ز�򗿴g�z:LrɄN�T4-�g �Z�\5z���$�0�:̅	(���P�+Ee����!���s�VK�����B#K��f4&���PԜB�#9�F���\��_ژ�y�������@2���t�Z�82;�Zin�*7o�P��:��j]Δ%t:ۗR�d>�x��A����j$TIt��7ސH���~���A� ���R\�fg��L7�ռ�q��V�VT���4[�~C�1P͑�M��6�@�[Q��Ø�˿W|�:��g�7��b�e<��ד���m�y�D]�=��e�z�#΍\L8|��p�p#���{�/��/�1���̱)�s�1L��:��.�������ɀ!JE�M&�"���''������q����Ci��I�xlxFe��Y�gΞQT�s�dp  ���m�3�����D^�P C���=J �D�͛�i�ti���p���Hf�� +46��t��V�s�@9'��\r�
z�	�sM�f"��͡�q^܇�|���>Ӧ�dڥ4��t�?w�ِ�v�Q�(e��Dt'��He5u���!k�I�eCgnZ"��3�V,m��m�ɕ�����N��K�qp��oZK"�L9�����!+��3�{���h�|�/.�ˠ�룖qg��c�2o�V�D@i�mF�o�2Y7�4�01�^����� R���m������fA�t �ZoXi�,:J�1`~Np�Èql0z�H*+��m��I���ι��7Ju��/z0��k8&�XR�:��?OĜk��w"�C�So��;k�՛a��~:��
(H�Co~%q#X�X�f �U�����f�{����+�ZQc�����N�DR�A4M��p���F�<;��H-)����Y����;�]�R)J�]�
���1T!8��vv�U.��Y�];v�[V��`�C�9���܎�۶���$`�Q7����'�7�j7���b~ ���#I�Ɋ/8i���Q����DՒ��N��y�٣��1�BH��,��p�Chlt\v=���٧Ti!�d�	�<�0��r襋�"�鴟GHr�2y5��+U�oWW���irѷp��7�f�w����Ȱm�>�,}�.d�Rٔ�FB��J������&@;7��A�[]Z��_���0�f`���H�o�`��� ��^Q0�l%�A�m~ѯe��Y%��a�>��[��J��K5�5=������D����-������X�f1�c̟ɚP��C�V�*M�>5��?�߭� ��&��,)@��E~,��9T9|��*����}\q��T-��}�����s��R8��ͼ �A`;��4"?Ǡz�O	��6֊�H�%$��o�������w�k��Ih֌(ja�(AQPո� ��3$H��iƖj�y�v�}{�[�ШM//��[W��ʚӚ��{�KlʟY����4�p��Hv�R6��Bk��)�k�D߭�Y���"�ߍ�4�f����വj�u"qY�M�0��ƒs�+ZͶ� g�D�ܰ_}�5- ��2�wM��D���"`�b�`��@I���^�C$����7�l^�EAy�E�}��   ��ݵk�6���@<�8&�Ʊq�Gr'ɔʻ��aL�� r� B�!�UE�Ϗu��e�3��{̡�ņa���?�e�>��\�p%Qc|3��<{�(���[&ڠwHD�1�<7΁���7A�}�&͎�t Q���>��AM'�=tz��x���D�%�����6d8'Flq?�"qSl8&�O)|?g��"�����d��pV�'J�o~����O��g��g��j����8�lP@&�B7/��D��Ά�	ť0�k��r�\TWw-*���Iu���κ�~����E0�u��#����z,���Ԃe}$k ��$)�c�tA��VV*n�F���#��(['�
�8YƆ�f��cT�u���ldr��Щ��t�}�[�H�6���1���p?��Z���$��@֧�e#]V[Y���X#ɯ�ɅQi��]��T���6,����\w�k��Ug�d��2aA^�47�����p�����A[�=cV�ڀ����0��sӈ���D��hw�[�D:�=� ��n�%#y�2'��x�xV��j�`1��m���<1�$��qml�&ln��/��\��$�"a+d �)5ޤ��m�m��ɚ��;Օ*��V�JZ&�g���w�uR�t@P�g�@ ��B ܬ߫��>�d�'�h4��:�h&�F�?����D����X4��l4�)��'��Z�T������.���2���/}�Q��
�t�z������ܕ�Wt��A��.�wx��g������SYeR���6�m���N;{朲�H��^�D���R��.��T"��H�|7��E���"{'A����>�r/�"J�G�>�sV��"�/f�Ά7���\��w�ϙv��1y9|�)^����Tf= a�oOۍ�$s�g�f���%hx�l/�Tٺn%ԍ�N�|D'�Gڹ�n2|���܏0k�U�>�kd� T0���ఆD ���T)�t��]�	QSf��D���=����H�CM���������L��K�� ~W"���6�X4X�~����=��8�=�����x�{ �����L$@����&�]o�T�h����n��~n�O}&9�t+�5�؁j#�U2���P��R@"Η�H�$�,AZ�_��+��S6�YcҾ��|p��:��%L���F?mE�^(׶�I�Yŏl�%�o"ĝ�b���JS���(�k�O��#��O���|�V��"�삃��ɨ)��t��$��@��u��!�JG#CcM�\��%i�|���B�QΏ?>!	�CwiL�i[�E9�����"%k�� D�\ +UM)S������ځ�4]HШBgs��h<��z�\_ww�����g���[w�!�
p�& ���"Z>"C�Z\��{L����r�D��u�ⶩ)-N"j^d:O�:eǏX۶mGD�<��֛���!uPJ���o|Cϗ�6�+`��F��
�r� vҷMm�]�3z�="^��a�%qB�ۻ��kZ�������u�f������>��''�hCJ��T<y�����Ŷ1�����5w���==<4lW�]Uy�#�WYd��(���OJi���>*$��0�H��a�� ,O9��4��v �>D�	��J �=]趙����Z�6o�s�-�$�MB��H�eTz��$�E6���r�a��wZ*��+��[6� rC��`��G.t"ce�h��Z	p���N��H9�#sA'4�I���b�n�שn��Uiɦ$"�E�f�f<�M5�ڒQ��2�����~7�AW�>�TQ`�������-_�mu��q�)�8�F?����C�tc���%C6���;��XO6l�/����0-d��Ļ�M)�G

�(�O��%jg�5XG`��!�Kgo"�g�o�Y���� 1u�$��D��-��xB�I1J����y �����- Hp*2{Y�=��sG����Xr[��N�^�}�떠��X�#֡D	�J��w�p���I��m	�v�d+��M�3U��%��to���t@f��́��;w�Id��c�Z�F�6L!��ًs���̐���6�߳�gf���AƑ�a�b�ؗ�76�浛��}6�]�v�vlߡ��`�Bu �� ������;�ɧ�'ӚJ3;���,�МI�u2t��������s�ĝZF��`z����;�v{ZM���VV��I9�Q�,��X*]����Ƙ������޿�~�훷�����Au�+Z�{�x�Ie�i�#�Q�T�]l����d�hDڕwG����h��d{��z��͹_��|��,�l��t4��sFE;��q��y�}?��^K����A�vi�"�&Y��*ua�}�E,�C�zz�'�d��xOgW��!#SQs' ��F����(D-�:'�B5�����ZIe����o����ɟ���]�6�&۶��Q��)'��-�tN3;���ǒ��u�<X�gp��eK�u�����^ZE7��k��S�����N�(����"70~�LZm���Wq��� �dx��?�,�Ƭm��N۱y�j�w�݅Z:<�bu!�ZᖑQl6�yӾ�K!���&�\�)*x4�������?D��i�`�a蘪&n]�9#�c��E����&�T�P��N�L�i������w���� C��( %����}۔�9��܊�7�դ��FDҽl�="[��AI�r.Y��S��1)���t��\���%D�y߰o����>Yܔt����1�o���p�T]����2J��A�ȽWv��m8�z��Xw�w������䔎���3�>uC0����!Cs/������p��}m���kF�5��D"6G|х(��us��9=�g�ch뙦��*��/������')pn���x���b��N���ƥh
M.M�R�`��.�^�s���r�� t^� �Xu {��I{��!=����ή��(E2�4�N,ζ���cԫ�Sgi� �>�ǝ^X����eo���ŲF>�2�r���(�M*S�TC�_bK��s�{Ϩ��l�V|O�\��6������^>�W��h봬�}��8��M �ZS�g/U)���+t���ɰ�|e #穬�GREׯِ�g~�7\����U�Ɇ���N7��&7����
^�Q��Hw�f�pRi�yQ�N�B��i�h3X�������E�C
�鄴#�4����@�q(�1j
J�AxF`.���q"]3������
]�L����Lb(���K}A���\f<�!�D�&�P���JE �e%��|�V�s�Y��Çڶ-[�V����U]�)w}ƽz�qY/�>�L2��Cݹ��V[
�Ȭ��� ��Yr���F�7~�3iŲw�wgN�mS�$�q��ɴ(�	4FP��� |���N�z��i!��bɓXߖ�H�$t��zhV�fCP�z����\\��G�UE�r3%6ۄl�Ŀ=���^ag���&�����g͒�k� 4.�P]s�7��w��Y��}�����7:t0�
*�{ü���8���(��9%-�����r�Pf~X���:{5�Ζ��5T��>霚ឲ���W�Y���|����'�[�YeŰ�����{19��U����2õj�;H�s�7k`O�V�������'&Fݟd$�U����a����M&��A%~��Q�_�H4<��[�^}�ذ��11���k �!��AP����́�ǀ��c�I^��Qy��|�SI��S��J+��z��r胶��9g��g�}z�.�.G{0�؎l&��.5�7��iw���ʥ�J�4 X�^��Z:�D� ��M*�nF��d�&�$2����scB�3�lʦs��Q����S�g���yE�?��r���9#z�� Y#�l�Si)�����t1gpJ�!ıc��DC��Պ�/9��"����8���J����(J�X�>'��&�����Q�`D��暩-۴x�Bn޼m�8p@Q�>��-n��x�׊�BSK�6y���FPt�A��<y�Q������[o�m켸�4���4���q/˚#]n���A�p��#�S��<qℌ��K,����h��;�w��o02��A,�uCH�~q�����:ۓdH��l��a]���X���aD�]$S���ѡ��O��Zx�)�F�E��R�8�""1e�g���0���z���MD\_Q�j�a< k���O��م@��G�1� ����]5;-�:Ǎy��PR�4Ɵ�R�=�>(ԕa#Þce&d���ɮ�Z��{��L��5�g�8v8�D=a?7�J��J�2IÛ�$��|�u�j��(�@4�{.74b��!��)5�!C	��ѴP"p����v l��R���'����(O�2H���F�*a" PZ��ZU�<j�~����Ml�22+F��qjE:�p�=�����m}����6c)wn%_'	�ƾ�u��$��qMZz��<���[�|���s4"�IcM �]��a�}��:dȎ��%��H�� �9Y^�+��F%�ND�c!H'���V��T����Ӱ ��f�j]�����F���/��V�Zӵ.ܡ�5O�+�5Y��cvh��;�-E~@RG�~w��g�U�j /:���4V�^^�壙��b3dՃo
�ܝ� uG%R��T	�cJ���V#�lS�W��u\ Ů�;lr�|J�VVc��`�x�p��U�k�O>�Lv����*5�A�)�
�C���P>���)���/���J�	�!x��t�ϝ��$:UO��,)[h�\��=|W́���;�������R��oF��ݲ�d둈:�z������u/������ƕ���\���dD>�U
Mb�dn�O{�O"��C��Eo�T����|h�T�G$2RO�8��LϞ�L ��K��<�+�.���a����+hҤ�9�k���$?耦�{|l®ݼ����������H�ZXѸ@��l�������F<��� 	�q��A�3L�a�ŉ��"2�]���v��k��@��ci
�����ի��?���B��!Z�hn��tN�YL
`ჸ�/e�ݾf��q�o�����ll`�ͮ�m�@<lv51�s	ӿ7�ҍz�J��Lb� �5��&5o|��O;�m���;��҂�;q;ػsʾ�g��˚/��-�n��A��r��5�����AS7��� 0�Ϙu<80"��[IE(ȼ���?�w�O�/׌;K[�������l�׹��tId���FS?�8[������2�]wAűc���$�=`����|�8
� ��pn��=����L��}S����B���p�����D��x1A����6�ɓ'�<���l��'�	�"�C��P\""E�W�C陨�EO��B��R��+ץi�y �0{晧#^Gp��<����Y��8�<��[7�z����੃�'�|B�I������z��d*1��kJ�H��8 �85�r͔P�9�A�v2�ܦ��鈆p���$���L�(ϳN ��RMA�f��$nI^���(L�?��ӵ(P����J:h����ⷾ%��:��tEj�
Jܑqo:"�-Ƒ�4hU2�\���dF��X��b��ȕ���Y� 2;�c�
�����42���;2��Cw��O6��Vn]��ʒ���� �������i|%i2m9&r@�߽<ֳ)�}�xR�%u?�+�D�L6�X�LN3n,�2k����Af;�<�;�D2g]#�Y 3������C~�2�=�Up�4����po�ͺ�]�yͺ<������"�*k����9���@k�Z ���-��L#x7] ���Pe�)u�g����,b�YI�5����w�hy�����~R�^��Q����Y#�6�Je�(�x�k�h��8�T)ϼ����} ��F4}y18�dV��|�)��������ʮ֭�0m�M�Z���\��T*#��Ow�W�.��avN!Ô�pu�[A��݈��8���~�d� qIZ��|�.�/�s~|JT$�g��Df��0>�:m3��;
��$(1t
�K�/���eo���)�id�h:����p����n�@h� v���+�T!��ZI�pnدtv�����������`w�|�	��.� �El�M��9b{�߫rs�q_R����}@�_�ꫯ��H5���߼���Qf�>a���pԡ�`Cɢq��._������s���F�8��׈����ufDG�-��А����^�/|f�b6q��Me���Z!���.\Ǝ:0�v Wʰ���wR���>��j��[����|c���gx�}�t�=�|�k�a��SD�U��u;������ܞ��� �Aܴ��+J|�V�(`��H�q��&�X���ϑP�v�G͂}~���a���wm�1��gz�Gv3�l��V[K|�t4�w3��3��	�Ŋ=��v���{��>�B�.YB�Y}C���biI�D]�
=״3��2����5��� ���Uw�}�ݖl��Q�칧��)�??%>"3&ɬ�0j��xM4��}�$}�4C'm�V�XY��Hp���JшM���Y=uw����!�H��1Sq������q֢ٚGG��ʰm��̘N���Xg��� !�MHW��e��`)�P�CD�F�c��21i����X��j cdr{}��q,�;�(نwXx��I��	�H�����E�>�Q��s�m~f>�v޻�:�y50O�ժ���=x�Am(�����I��x*�'+�?��?��9����&;s�s}/�S�y�j���?����K���#jesOG�����#W�{��=�����̝ ������}�WJ������jذ}]}6�ɸc��ɼg�	��epxP%�Ϸ8X.�3A_��:��[�He���Fd���ڊ�-,I��]��\11�atxH�t
���n��5�i%�Kjͥ���)c$X��]������Ԭ���t��Y+}F��ޞ.e�0��&i�%��87 n&j�J&�O�&W�h�x~���{y���[�H�����^���T��x/�����{gh���{��H֭Tw����*�Wș-�إ����md�N���������7�Xw>��{$�q��m3]9��_��DV�<��+�>.K�$�v�8eQfLY)��F�!�+��F"]OZG*gUGH��5[j�X�Ј5�9��lѬ 韔b�~�q�K;�-Yqf�F{
62���I��[	[�@���O�D�~_�P�1k8�L��5N�����0k[�z�S^�ޮ��_�r]Z�C#(	RWפ��71d7<���0g�>K�UCfu�R�T!�1g�����s�����Zt�Zo:���~>��5���z�̊��d Zz���d2j4QW��gWG>�i}PA��y�^}��v��;8l��jd%��P�
�5���#�l��Ne�(3���w�}ʑE��&q>�ޑ��,ϳ0;X�1���'�Պ�'�<�̟y��X�S��/���+,���Vt��l�_��c( qK���'v�������V-<��&���'��$nɞ1If�Z�j�F�)�Wہ�x�`H�LfS�+a������-��ҵ�63?��F|NτF?�}_�/���	�&��q\�"{��޼���\�f�/�����Q���W�ط~��ʪN��рJ��}V@{ŵ�M��={������|Ʈ�l�6��~�kM[XY��c��x�~~��&t�d�oܿ��1{��cҁ�Q#`6+;~`����q�T)$��7���Ɵ�A[�{��RԳ־Xs_�:]Bu�С�̂�®B�)9�7���� �þF˔����<t`�ﯬ�� b��Њ�w��3��7o�	�����ш����,({��_^���8,���Z��S�U<{������t7����x A����Q��ᰗjatcwO��]��w��M�s�V�z'��RI��S�k!�ތ��͚�\p}�W�5s�`��m��l�b��Wm����Q]�C(S~M�h[�=�����(���H�vG�e
�7�(3*y4����[�s��57��p�¦�muPD��1wiҵQ'lRݚ�vyA��t��=���c���a:IKH]���5���3��QO ק�]=�2]誮���\_oT"&���$�#/�.�c��s.[vn�a��p[��h$�nl(��h��/2p��[�c����.&�b@H�s\6�u!?��I� #zՍC����s�+[&�j7P����#�0�A�c��6�����7j�̹��iTȱO���==m�z���y������#G�yw����I ",^�+\aԞfI'm����g�.B2��cǎ��NWt(�l�������F�u��R����� 4�B�dH�A�ρ�i���}̂����K�LJY[�9wwv�|�1���n�cn�ds�4��RD0ǀj}����'�@<.kk�Ō���ۘ߈דw���޲�yDFZE�Yowi����8(��h�D�'�nXJ��|��1�Œ���	z笴Z�aӳ3v�Ԩ���^��.{�W�ڻ���G��k��-A�_�;M���������Oϟ�?���+�}`K7@y��M���|]���|�ܳ�Z�e�H'�S�>ԙ�������+�z������e��`������\?���C;�AH��n)i���a�F��n�g	x���I���J��&���������;��4\�q�R�2t�k6�@�ԥ3�w��Җ+h����#Zz�����wH�Vc�.�B'#��9�P���O��u�N;u����W����5�B�tP��ʈ�{��2*u{��'l�褃�4��V���]$�>�l�r{���W����^\p��l���VJ��!~c3�G"����X���ʺel�ݱ�^��7D�������͏mzyUӪ*�*�^3k�;�A���ݷ��z�Y�#������;lmN*A����S���������vZ��Q+HL!�=YW�)Ѕ���$A3��m��C&!��E�ɯ���̹s�JwGA=t2~ <h7�)8�|؅�z�f炮�O>�y������H7/i?��2�d�Z|߆�D�l	��@�Y4� �{��I��j����m�K%�Dk��p5j�=	��^��cϣ5{�}���_�?�D `n��_~Y>���}d�42����E�V��>u����tҏA6����/�S�]���O=$c������g��=������ZD�a ͥq'��s�ȴ��l#��ܭ�����nSխ�p	�n�a�'��s�u��6����d*L5�s��"Y����&�H����.�Z�ʆv���-�F	Z@�Gb�7���}�������3�̬�̍|z�dhID��_�8�$�b<"����� �sS��݉.����پ����G��1~��%�x����U5|��"{����f�ST��ܚ��õ�[6���Kjp	��G7_֓�'������,�/�(��Za㫕:"L"�����-X�����-�jؚU�P�~Yt��B�qY�)}-k��t�!a^���݌I*H��t���OT����	���P������	���
��tq�t��X|�H�P�Իr��	�gZ�$���a�TC�)x���߯� �ri�jj#pdN t���,�^n����b@=������# ��5� � >��	�駞�y��W\�.qʭar�!J� B�W�%��e�1%P��w������"����GߓT� F��{(QoټY�Q�e��WJK*�SZ�޾��ka4��,��yγ�s - 2�i0[��NCMKqc
7�ڍ��2�z�n��)/k�Dݠ�?G4:�� ��JOG]���Rk��͹p��nlʈl�9�qMG����2rh1���$rL��Gw<��pjݍne,(?r�ȼط?4��ZPw����;g���JJ���&�Κ6��0.���b=��NK�:��q �e��O_��&U[��vLٓ���R�a��;�Rf�'?����ЕK��G: -���?j�qp�����h_��#������`ğ���	���d[���pۺY&-�\!%P�P��UB�|���y������._8�Q�v��A�)u'���IZ<Ť%A��vtR�${ �bVt]%me��@F�d粥�=��3�{�x�:�^d�Ut��sf�����WOnxlЯ����>e���go������#n~�w�i��:���`x�O�6c��h�y�0?m;ǆ�mZ^��G��p�=��~����Ҋ��:P*7��:g#HA�����/���u��� ��S���6[�u�m�ւݿ�>)Hܷu�^y�M{���R9��bJg��8�4�d������Q^�s}����Tn�/���#��c�n�����y�9�c�O�f���ߋ][��#Y&�����ò�X�4�B�?L%g�##n3����S۷���w��. !;O���e�n���1=&~uG���\�z�ۍ ���R�P���Z�T�C�G/�1�c��C�! E���	�Ltb��~1i#��k���.ӉZ����'��QƥQQ`�7J�r�*(�u�,�[�@Byz��/(E�G��> il�M��̀bt �U%P����t���d�2`��'��u��$R�U3Nw(����(v��s�iȁSοy�1�8�z��E�[�ح陠帴���	��
�����w���,��^�rY�w9��%#�	�k<�t~�I�-$�"e�ۃP�.E�ӧ?W�CHH�Jр���n퓋������۲߫�:l��&= .;`�D��u�RC��,4��yK�z�+�e��?��F!�A�������~�\~��~
�sA��&/YU�N=�L�Y��CTV��td#a�Fm��d"�hQGC"�� '��C�疤��G���~�v�p_�ۂ�U���]��4��t��ݲ�U=����Տg���15c����.;R�D�e�8{vm�'?�Ʒf�e+������ᑀō���2�18e�Ƣ�8^n~�x���E�$�^8jn.�D�|8�dD8ڙ;�:�哉��q��	 �F�ߤćT�����T N륢�G e``H%U�I�Y8���2|cX ��\.��7����	$�aJB�I[_C�1"�F��������w�� t0D��3�ȴ��1hd�Ȑa�X(�X2 d�R��a!�Լ}���D�O>��/F6�8dl�`\smq�P�⠌���o���i=��s�S��}o�k�N)4Ϊ�Zk�U~�����^���9�D�`K�:&��y$��ϟQ��Hʘj%�Q�7�V$MDW$�Z6�9�a|f�N��Bd��!Tn >��3e�D�;i�xh��d��&ӭ��|Ϛ�c4��x��"J�X��>�����/
����q�Ú��Kk�^k7I)S�N���CK�>QTS͊�L�v��m��V�����y}���^wگ��륧�ry���]LG�꒻~��?�~�ʦ�/�����q�� gj��Қ�E';����,<%e���Q��_8��ۍ������_���7���_��SK'r� ��J�)q�[���v�����":�=�@�&�g�-�M��o�w{�:��Zd��}�Tk%M�јQ�|���,ء�ۭ�������n�~��wj\__�-�u��ZK�Ȕ�U�C��7Ɲ�s�ŹEq��+��ˁ�~�%���߶0}ˆ|�nʳӶ�Ȏ�ڼ��n:ߋ���:V��|�q�z�V--Z�����	{���w|=�����LMˠ��[���3���쵾|6O�t[�d�ZEzqY8��0����6?��\�:rIM�Y��^3��
Yt�Q�e_�cSY<�z��{h��i9)ߓl(©2�Ii/Eݬ%��g;֕#����|7Y.�m��X\�=Ρ��t!;���%{B�aPihZ��1�٨���:��fhL�q'6�� �giJ!��|у���?;w��8d�۶m���	{�}��[Ӳ���� ������~L@�4��n�B�����W�|u�O� ��㶧�]t0�y�vВ���kژ����{T��9�p?>q�&��e����.q��dn���Y��a��*I3�+���n�V�w� ��!`�:Y8|6ׇǏ���1ӏ+�c���=��K�q >0�/�Z�����>����_��^��z�ͺ��;�C�O�v�P�GL�ɭ�;�H,�"�u�� {l=���>P۹3��Ibq=���d?�q�����x_2��ŋ�O6�V�J3L($j�q��S� �T_j���.C�0�LDMt������oW�$�����u���r���z��v�Q�[���ʿg�|�-� ��P��:!h�������47$ qP@'�2�F��0�_8Hkv�������DR^���qY�,,ng�\6BG��RC�5t'�J�OV�1p<9[dp|��X��?�[lP�G3�����	i.��D~��f&��'�d`9N�!�� �T\�D��]�)�����r(�<������u��o�	����L��r΁����	ta������IN�:�44���{�h����2z�\����C#��H��:$��&�9|t�Ѭ�{�HXh�=��"Z�M�{Ùs.�2[���0�p.!cȘ�0����?�����|��~]S��z8. �/F����>���č=�G����#	��� ���8SA_0�PJk��*����DG��l��"��8
���ϋ�`�4��Bl��#<��r<V���I���Z����Fo�@"��Q)^�r!�Бy9͝n4���ޤg�qG'J�_��)+"ZE.�J��6�͵�@Q��I�Q
"%�Iw�/\���>�:>d�g.	(l�)8h(��ّ��.5NА W6)A��3���V}��
F��"F�2w�vm��?�O�؞v�q��%9�>ی
̒���X,��9'RN3��h-=��?���ٿ��'�z%��Ѣ�	�e%�+o�ĭQpj,q����f%߫K4�uv�D.��2����Q���l}��~�5^L�I1Y���\�8�3�˲I߻�w������{uƎo9(�rJ��i2ȸc���?:2i+KE�9`���@V�#mK�M[�ۄ������W����>
����ڈ_���#J�D����z�%����|OgX[�����*������O��*~��SM����Qe}:�}�����yޖ��;���*��}�Oߺ���/B:��$�EG�_g]�Ye���1S4BI�'��b�^�)*�eD����QU(/MC�\�T�::�b�w�J�s�z��V��iC�5Ѿ	�����m��}�F��p6��~cj@!�+� �/7����F��p��l����<,Ё�����ő	#�G��2��k7�'Ț��M�!&�q���H>��3S¢�Pbf@2^-[p��Y�����wn�x��%{�n�N�A�;/��?���@=%|�$��ؼ�;3*����wm�d{74X���CC�D@�0�>#����$5�5 z�<���]�הM��m��`�2'@{���}�ܱ�T��|q\�$Y&pɡ���H �).^��2q=J$u���9d�ϗ��*�[���6?�b��G�!hla�+H����$B�7� 	������y�/�gL���a��'<3�!��R�Ik�Hb��b�$g��~"�F�m�T����3��bh���y�W�ɯ��~� �y��TK�V/$�����I��6��򠻿�A����e��d�}`���*4 �B�-��f�D$��"�L�ΆM�	%��iL^T��7LG��`�ˌ[��3S�����,n��GELr��]�h�^*���M�g#��B�k^�Jn49/&|�y�	-4�@(H��H<r-n�a���<峀PD8CcOºr�J=nwz�3V4&��&e[�	H��L�:����	#t��)���&I����_ڄ�C�e�B#NJ�E1l�˧�<5�����|1��"c�wqm�|��w��m��G�s� ʽ�:y�Q-��Tm70%�l������a8����9�f���R4���>"/�� =2����z{�Y�ЉJ@������$�MFt��]:' ����	���W�jG�H��);�Q[Ֆ��v�?��]�;�)WЦ�~ ̤��-��ESӲ����ʵ�[iDݘd���� <�C��Aܹ���H<6t|��5�ϟyAܖP"��J�����Gy�z�;�PE�zZδKkUA<�F����F"�i�E���Nȥ���}_t<��}3�@���hi�q�-?ڍ�8w8�)��LLiV��w��:��(k��ǜ���K���C��`��AO9a�#������v�6mWn^����:�k�*����Uw �������7���l*:�zJ�L�ݿ��J2ؓH�&�[zykT$fnY��Jgz�6����+�u�'�|J���}sn�/^�b�/]t�_��z��C�x�D��qMv��ȴ'^�o�/���j��'���'���Zh`M.-���^��S6�t�ہd�d�b��m�� �U��Jr����mۦQ�����p�6���q?���y�a��}�q��I�&!�Bك���o<����wT�O4S��2hX'eq&���x��'�#:�:�["~ډ����(镦ux`�B�q:D�F'F$�&J�9�a�sZ"�q ���\W�uo����D���ߝF�Ҍ�z���q�O��hb��)D_��h��18����w�y�#�>t{����TtkJS�۵�ʤ|_�6A#�罴�`}=p��Q�c@A�;���<�Ur�>� �跾2���%�J� �H7��%�@@�M�����/|m��|~�~�r���O�YdO�KG�������?�
��x�	;u�04A��m�h.} ������ފ8wy]�<����x�1@Y�Ƚ���H�����V��������C�)U��ԧ���yPuCw\�D�|e�*5�^������@D��e��m*�:�'2)F%u?�QppIW�8���x��Ow�z1d�o���a�A�?��G�mJ:�ӑ�;��`�^�N�L^Z��s�j%�)|~�� >����۹�(����"��T�ܾ����ʎ���W,����cA#z��l#�:������%�I���Q[�3g5݁n�]��-�6��a�
��kl���2e���a^q�_曉�.�U��=�Z"�bҍ����ܺź�	��J�S��J�:�1,�0n��Q"�%���28�P�_\4N��8w��6 ���&��U��^kD 0�q�)"��C�&t d�."^�W����JK�EK2�?��	�/J2��ŝq�J�!�a�Q���0!���H(eP �}ǄQ��η�v�y�a�1Dr}����D�X!��gl2�+����� �C�u�P)�{2z�x��+W���!lF1
�(%S��܃�E97"3�=��~@>q⤴ )٢� �d^1VG4��Ȝ­l�R9lv�$"s:�`��u��_�g��L&R���>���B�ƽ�Zc�sLs<�I2n�� r*�L�:p�ÛF̘������F:� �����QK.����Bt��w�tb�r5&��pަ�H#�D�OZ|8�F�������x�tdp��8�ꦔ�	���8�ͦ$V��5�ԟ�f@3��������.$۝�l��G�:x��Pp����9�o�z�ܲŲLY)/K���w��Ͽ�������Egq�\���g/<��-KA����	[w�],�[�Z)D��ƅ�D4Q���ɖ�U�3~>��g�:�re�ܾw�x`��,8خ-�ө�i�U���~i���֝ێ�+v��E�������������?��A���6ߏ㓛$[��rpS�^+�o�������e��dT����œ�٢�����=��75�-�6�}�O^~�Z=��k�v]Oڇ�2�o~v������|�V(i;@�^���?;���Ծ�Y��J�f�ʚ���{���6��*Q4���;��Y���}��Sv����X��9�H�DNy`!L�2E�o4e����
��#���O>f�rP�H֨��D��DN���'�p���L�S$��z��8`q���xܙ|K�#��d�2��~m���{��|x�c[$��&~L9@��JC`_6�{d��g!�448� ��=���o=����y;��)?�uQ\��9ߞ�q�xA�ؾc��&* ��0��ڍ˾���o�iF@b����)��D2cO�s���/����������ߨD[��9����v�c�����k���!T�<�jS<���W^���6�i)d;	�nD�) �Lm�`f����ݻe_ ��CUi��ty�TQE�u`Jcý{�0�	�o"���5
`�����3������ ������9��ɧ�>�� ªﱞ�����\6�i���¬���\�*\N�9�� `#рD���e5|�@��X�Kf���M2�2q�t���R4����O
����45&4��'�����U*y��XQ�V�we�$t�oAb��c�{��6`r�������y��l�b����W��!�������/no�2{���_t𖱊��jLUx��|2��56݁�a�w#i�e�����=�5�BU�I��z��I&ڨ?���(֪�"�Z�+��V��Fh7'��M������ᛃl����Q���+�!!�\,���H'��.g2I�!�� ��΢$K/��<
�56E�y(`��V��JQ�;ٴ N�l&�G� '�@�M�FSp�4x��N9pA�-���(�Mj�T��}�C���k��(�^��/@���sq@|D�=i~O��f5�8��������t�|B@8q��D����2Ttxc�dt|�1&�/j��gG3���0t�L5?Ձ����d]�x)�S�1q|�gĵ�u����15C����L�L���}FΟ�z4�p>��t�3]�VZ!��f �5�UUN��q|٨y�������qN�U*�S6����J��(�ƌ�:z�D����]���_5}&ݡk�yh'��2
aP|-�D7J�Q����֬"���xT���F(i6�N��!�dT�*8|2BD�8�đ�}Kk��	�NW)t���`�ͷ޳R�`i����B�������|M��7Һ�»i�zޝ)�:����d{�\L�	��{��!��f��d2��u���Z��`=	wzKs�ٛW�kvq�~��v��i��4f��������d�������|�����y�q�]���s�
�19R�NWK��ෙ��g�/Y�kкF'm�I"颤&z���+7�~�g�&�:�j�CZ��޻�~{��7�\k` [2N�l>q��+�E�-�p��	0����C��o[o�˶�I�5BY�{1�k���m"d��� �٧��C�vX}}�ڮ�7�W��s�B �����{ڝ�D��>��M�?%����,ί[�%�x��g�Z a�4���k�uI��H�sY�_� �A[����r��t�X�,Wܾ@�����d����c�X# $q���+�?����!�IN�yh1}��
��6ubbRe˫W������0���踪7T��c�swdoI�"�ߩmS:́�^^Ui[�%[���k�y� ���aЃd���/�B��}N�����\:�T^�K�|l˓O?-��yQ��g$<���S>*�.c�;8o|'
��7��N�d Y @�9�k�}�t}uh���vil	i�1�F���z��!�ǌdD���3�q5���C��@������a~v��m��8��=��@��y\L�!4 ����uF����^��=�B��g���*�=D����M<��)׼Oc]�!{�M��RO��b���`8$o:u��N����<c?�O�O�9P]��N)�'#��/�������`ZѴ��&U��)5!þ��'�L�SP 	� Nr>~�� E���L#�Z�1��=hsj$`C�\R\�xJK�jZN�V[�$��h��Z)9���D7*tWKU-�lԴ���`�Q���A�D���E�=�P'J�����`���#��/p��B=�%�4ʣl$���zhL�����cIM<�����N���i=h5�$[myn,�����}��-2V#6G<]�fh��`��R��V�"�� �\�>gCa  m����ݣ�a��٫�S��D|�G�W���ں1��c1Ph)J�ǙC��ޗ_~�?��J&\�ǂ�shk�����ԈA�(�p~̮Zg{JFo������?���>��3�fCf�S�P�}���䩈X�}{�W�߯�Z��Kw���TɃc�8��G��4������@�����
$�΃��������J�C�X�P�8P�FFe@x��e��=.ŗ�5�H��Ϟ	����p�"9��آ��pdw��)>%�����T�-�'���BGֶ{477{G
 $�����2T7�0e�9�5�MMf��Y�>۲�{63�<���t��K ڜ�*s��n���%e�g�V���z���s[���Rp`RYTpsd�[�	�m��N.ow�^�:^�������������D��d<Z-�o��$8�ޚ���߽����tݞ:��U��^qgXEnρH=�Tg)SKr�B�L��LZ�n�kO�e� � $x�0Ć}]--ݶ�M�̆�Rsc=�U��,W\�+Xʿ7Sp��HZ.�ike����k��s�X/ۺ�*l��{��O!���F&�m4���Ų��2~~$K���X���N8�x孷��<�F�S:���	6����/�9%ԥX)�����lz�m�;��?G�cR���K�z���i���%�~�)[��J������Ųu�Q����o�����^)�-Esv5�]M��^&7��[iU��EVʟwu}����U?��jY"�������-h���J���K��K�j�_ϐ����6��u]�\�F��U���c���(��@Gso�A�Z�KҼr��L�{	 @�T,j�
v�c�H�Jl��w�}v���m����S���+|�٣r��N�o�g� K-�����q��49�!+Ğ�n��"�!>��
��M���}�wmttB16��!Ǖ	��?�c��ѯ�3��ok�����8����;zT��|�=L"��.�����v���q�?u�� ~q�⃎��J�t;G���u�?��)-*�Y�L���p����	�s���, R�9>�r0 ��%?�&���h��d5A�$W�3�;8���n����9�J�We���h'�b�E��W��s��[�gH�̈́f����=5�H�l٦u87?��P%(�9����0*.?��zdp�u����� �1�h���f�HM�uB����k�~���
ɦ�s�#TN�f�7�
���8���3
�hP��o (V��G\ܟ�����?{�md��u�˺oP*���RT�(&���	��<��������1S֞�Ҭ���bMh��uM3)���"ߨ��<⬕V��+kJ��0���z������.�`6*	�e���8H��x������{��xW���e2:?΢��B㈗���lI��0r\�Kw��Q�雊�f�fȝ��4�$�,�3��N�>'N���@O�t��X[^���L4�>����o�>LzK�0H7���<�]�w�&w�?����gc�ɸ����UE�|SJ�yJ�6>�`X��|���8�=}!���hI<���!QY�(�c8�nݮ#���q�)"���B���$��?�ۿm����=��{�&Bނ����4���FϜj���T��q�2R��Q����|fg��M�U��Ueq�o �}^��1�[��3�P�}��?$?%  ��IDATsPݠv��eC��QM���`���pc\�!�%&Ν(�c1��sJ���< �Bg&%8�d��w=ʰ�`_q���8ƍ�q(#Y�f��@^ţ�s�Hǎ{(��f��Y_q��Ͼ��ߪ~��:IFЁR�Rѿ'� �PU�'C�I*���+|T��ݰ.:��Kd�00��rM�N[��������Y'#(=x���'������mV˚�,��Y7�ZeH�$���̴I�ɠ+�L�G��|�m����Y�p���z�;�c3k�tΏ������e�a3�8�/_�F��N�d���i˾&V=��N�R��Q3��rU%��M�g��!�̓�,�sϵ��<Oґ�&��$<�sgp:�o�ν���M�:}���T����U�Jխ�vll��6c31$MG�љ��{�������o�*�@g������w�g���g�;��d�3��O��~`�]�98x�w�M��ƶ����SRBh��5R�&�L�;�����o����t��KBU"�(.Ή^�p��[��{�N\�Ҋ��͞�w[ i�����z`�́���	��%M�i��e�myi(͘5^A��)� {3��!�V5f�;��T�{uaZ�>���!i�xF�>�������\-�&�r�y��9O�R���k^�hN|=�5��'�"Ԉ�5ґTLLC���ISG���s}�M׻]:�h��|�ځ�D���}zzV�ri&����&��?����?�G�	��5�\��/l0���zS�-���R��~�ᇥ�8���?o�ƤN�\@�_�����D�C�%ӘIV�{��/U�X��D�?qm-��~��0 �L��Ir��%�"�֋/�`�f���Z$��[���c}Q���b�^d�9|�r��m�EF�Rzo��Y�W^}E����o��'{��㘲��U�"vOs��uiZ�{L#�8������]�g�Uyʃ7hj�g/ ��6ሥ�t�됔 @�2��:��(:�k�tc��Fr2�p3y��c�8�1�*^�����n���|?�'��Yvw��jIs���o��5��f���zK�p���/�~�=~�j|	SG���� �w��R��3�j�wm��<Q$��Y���̂�=yb{v�l��\���+����+MTWJE�a�Qb�T�x�㓠j$2�8�����D #e#��3��s�^B䦑j� 7 �ㆇԲJz���b�$�r�h]�А�$�@�ql�f	�J+���������h�T�nF�Дg��������T<H���Di8�P2=������ �a �
2�d� tAg2�$9gZ����o>,b1�CA��	���o��;~\����0c\ؠ��:YS���3�u�)Q�� l2��<��mK��5���  ��N.�JJ@�=���\jH�D�pV�̥���5�Q���d]8x�F�>\�h��y��:9��ꥠi�Le���&<~γ�OCYJ#5���{�J[$���q�4PpV˫����C8Y��d���F��r���u��u��G��qz?!�Q*-��oQG��� �d�yΚ��ڢ3 1.�]vԡ!	�E5f!������þO�S��8o�N����#VY���֜m�sssj�� YTdґG�~�[�0�x4�9��JD�XU��GN�����
� �
�8k����V|� �����Wh�F��#��`��R��2�;e������&��e����L�hd��1M y��jl�bZڐXY��gOk}[ݙ�d�j�<?iC����|����vڝx{ã�&������7��Z��Y���YJ�Zr��N�v$l]I:����Y+��F)?CfQ�|w��R�ЭZ[XQ���˕�DyG�N���8�22`J�¨L4�?�C�9��|w;h����]s�U��ɥ�����[7��w�nC}�~�3έ��ȼW�d�(Yҟ}��}�Q����&���s��T�gߚIڵWl�Nw4�z9�_vTd$�
��פ�Y�G�Ih���ep��6����3���濷���AHX:�~��]M�As�Ӓ�"�M����ي��8�<���b͐��fqV��r���]#?��a�/�o� �(^��U%����%�^�&�Lϭϒ�>V�,,,*�#��D+��p������ַ���>}|��o��5m�f7�U��A�HQ3�&�����c*?�&`� �;�׉=�ч�/\B>�ՅJ`��r�۬v䯹�ZufW�AC��>G�Ʌ��_D��JI�,�]���x ��y�u�鳰ǀ�Q�N9ytt��	<(Ot�o�~�>@���C�)�j]Pe�f�P�>ėp]��c*�;���kПD�r�W�&'/������| ��\>4���u�ܖhF3���IP@s�5��&D������eQ����ޮ�hP�W����1�@=;3k���H�0%J5�� &D�x�MD�sp��̶��&rN��>OE�6Q�ލ�8�d�ͩ�9�>�~���P�ת�Lᙈ�g��|QJQ�7԰�;��c�$s0u����Qq�7�۸ÇŎ3�r������R��l�28�ͨ$I���|C���F|�d"��#��*� ~0�)�G[b��L�O���^^YZ��A����s���C�q�;�`4��a�|��Aᢐ>������.ifq�޹�J�{�^"�;�A� �5�X��o�C|6h�� 5G��q��X�s&��p�U$�ueMh8�		���ۻW��X�i��:~�n�Z貥��u����(��	O����=��_��������m=��C��FY?�g�H�BN��r����x��EѺ���<�ŋ�"F De�=��z�.�wcM �HJʐ�[[3Q@��2�%E����ġb�p_h���-pf$�[
YL�Q$=�n1y$L���dTg�c �R	Ϙ}Z�$���x�w�1�p�j�~�s�kl��Fש:"��5��.Gޕ���y�?����It+S��h�K�� txD��#P���W�Sb�kV���|-a%w�K�+j���iMf���3��9���u_w�e4�T�����n���v�o��S����� g3�H��7:�r����nw�M�Շ=�ɣ?������կٟ��Wlhd�dC:[y�K��{�K���]�g9�{y�P���/�,�wln֎N�s���gJ�6��&�dMP�Z�^Җ)��qYq���{�l̈́�����u��N/��Y��*��@���$�g��d0�
�'^/�7��e9������ u��je�Ȁ1b��>b#���䭺���hW6��qr(��f��P��XG[������k�����?����W�c��g���M���RH�&R��^:�n����I̤�?���L����� f�*BF���46�B)�mQ{�]ϕׂ���������\hH�~�� !�^_� ���g��2,-/�s����h0DCI�F�wup�3$c�EV�����%�Mf�T<�3F&4d�� ��y��i�XJ����L��G��������l��<*&TQ����4��haoO� S��A�w��/\��j��r���h��HJ���	�Z���i.�Z�f������ڪl�|v1�BV�J�,>~"�%��=��Z?���>׬�x��h��ᾓk�f�Sxv|k!}^�|��ד߁��f��(��А2ᚹ	��];��xF�m.�T�8���iZ�O��k�U���5��PZ��e|.��@7K���$�R�����x����n�I�� �������(�-���/֚,.<w�����{I��F�ꬦ�����%!�4}'*AG�ܦ��i�t������b��Ε+�T���Wį4ID�­-����K3+~Hf����
S7r-�����It��aBP�DT�H������L���
@Q�v=�8�(�k�Ab���"��F�hkK�����������f����B���H�%����O��
�[��)�V*������FZn�q�&���V����������K���d��Y�׫�'l��R����w�7��k�M|�S��(Y�qw��AuS���|�7>e~�~�a7��8}`��X+2�8�8�f��=��c��y�95��<9�@脈�\#Q��߭GEDzG�qSL�iI$�� �����$��gRVg���.�5��s��r�ͷRU6�k�Ӛ��]�{��O�1��뮽N��D����~�Am��/���"d�����3�9�N X���Z���~��� � G��G��S0�:��v��Ad�Ec�0X�9"m�Q쒃'"h�[�EM���{)�ĝ�4�(���������x�4�i�` �/���%E���u���b"�r�EqunDn��7�Qc<�ș�^p�q)��rF�m�:��2Ī���3�6���;Q2:�k��t7ׂvA#T���IJ^m܁6Ȣ1�	�K��"�-6��l�y2�������Zjfl���C�)+�!O�}�fSy�����6;1�.ӄ� *�8x�H�P�:)��-��V�1�{�^q���y{��OY�����߆�P�H���)��B�Νo!�PW����V+d������l�[�����L�>玺ǆ{}M��ꀼ���y[]����[^X�Ƣ��t�m�%����������nߚ�ʋ9��}͊��"�Ռƪ���UQc_����/.�P\9үy�8�*�IB��{��۟�-�G%�Ξ��=Vw�	'+�()��f����E�ɤ�� ��|�Ə�iC�Z�>K+s~��I�쑙c�%q�$[�lD��!�@m����2+���1�1���D�v5R \�o��1�4�)��>,���${��qM9�G�Ab��
���[�<��[��IӖs�b�0����s�|�\�ޣ�84		`	�����Ç�Lz�1�	-��Zim-�.�R��9v���� �������]q��޼�V��o}���ܳϹ����[�Rć>�!5R0�dmeu]�� �7�P��ƾ�ʃ��Y3��8�I�� �T�}�U�/6�FǍ�F�� ��VQ3	l;v�j���^�u� :ũa^�����F�p_�3�\��1�� :2v��y�0�7{��c�^w���p #Q��f3��~_߀��ٯ\K�@2��7�i��[�|��ϟҙ��oSQ�U9]��#�=Cfu��u7\���c����aCӑ����a\a]C)��m��cf_H+rhH��g�8��K��\��ilx�K�{	���.�Z���,$��]����# S"��.�G"��c7¿�D#y���L�*s��ik����s=;9m�}]≯Bы*��@���Z����Bg�P"͌��H��$Jk��_� "�}��ସCTx�̴8]���|3�Q5��Б�|1��!6��p2�8Z���Mը}_e>w,iu�z:�$F��#tS�� R1�!i� 2�,J3�nz��>����7<i�MI�!��&8~��-"&�+���_u��]�	?@�ش7�|�:¸N�Ā��Ò�a�q<��-�6��^x��p֋��G�n8"Y��S"��Z�=�@��d���&�(i��(�q�?ƅ,��y��ub�-܌~�� �´��s�� mDd�6u�S'( Rr4a  ��"=�^a���h���}�S~��.���2k��{��k�hDp<�mๆn�:���@P#����@���9E�?��g=��Cc�D�"dse)��eh�����#\γ�}dx�q�;��Q�V\�r��0"�����#�u¸�x�L�'�n*h���sң(P�*����I��5� r����uj��H��Jy	�&`�q
pW��`0A����{k�B)0���6���J�^��̶����cK%����� ��ƪ��fE�p5T�E�5T�4��Ӕ��9Uq0�'1��6�;�\���%w�k�A������97��;�C���=�g�e7����{ﲭ�mdh�V4! �1����dhZq{�q��>���H�f�+o��ܴ��P]� �����v�;;5�Ҭ�Qk[u���i���v����ց<�����;w颽�	�gG_�uz���jq΃�FZ�:;4M%�H?�K�G2�����*�&K��$�!SC:����ˁXY��񛥊�\��4W<(��||2Ҏf&��ԥ)�֒� >����YK5�z��.kzj��Xo��oJ�	�����vp�&{`��<�EB����6"�PԼ�9jD��$��Yi�J�����6���ǣ��Q�P�T��"�@�|fnhk]��P*�vvv֕���� q��3��R�8���"k�P>����EA&@�3F�u��~Cv����0u���n�ю;��FY?=����u
�3ܧ��uw)0%�������`���~��9�����O�'ـ��T�y���7�ѡ��g|�ӟѸ���zZ{��`Yw�=G6�p��ʥ$H�<���;4ݠ�Q�h���h:�ARg���Q�����cKٙR�9�;$z�:�+���`;�rIFp�۶o���y�P�x�4�`#H4q�|�� i6�=��
}��
����Ơ��=�h�)�y�,d���� �(�jX��e��?�v������h���S�y�)X���f�^�_��DI%c�Э ��}�+�Q����VqI�g�
F �kl&mxt��$f��.-���x�}@1ƋCv��	E(Yؑ80��/݌�P��D|D�	7"�^ii7�k�5��x���s�"ku����h�����S&�:��E�ɐ��)����)�yg"NJ,��f'�C�At$��0i{��5�vR*i�}�^�hF���@������4�"�2�	�e�&͇&u=?���8�ÙLf��ƃfS_w���������s�Cw�`�N��`8�K=�y�")�x.\���_�n y�Ώ���ac���sfl�:�<�}�������7�l{�|(d�<�%�$�������ȑ�@9�r9�BW����ơ 2�żљ��=�ܳi��q-�'���a̘Z��'M����
�n`)3(y^H�`�y�uם�y�����0@��RF�qE�GA�2�������d!q|pA�D%b�������Q��p�?�~ݱ�σ����+�R������yL��� �c]F@&���'��l$��������i���I�����M2W!)�[ �;���Q�%<®�X�n�Ҋ�l�*�Pܐ�YQ���Jе:�25�t�w9 �l�Y����4͔#�y��j�H��������Y]x(��VY���K�{��;�RE]�UtS��-I�ZX������-/Q�\��Q}��KZo��d�E���`������k�l��kli�l-�};m�E��ϫ��3�f�����R���H;h��i�����c���|�}���$˳�6d�R�r��z`���1`GN���Z]]��wv�XGw��V�d�2���(���0oiP'pL8M����埦���4c�5ӣB����^ye[Q�h4�5��K���w����S\U�mɿ��� �_�R5�7=-R~�OFSn�TUc��Ң:tD�j��ak�l�f�.�D"𬱃��lգ)Z��~�},���,��O�K�%���mA�)!��˙�Gɺ�"��H���r4���|]��**�{p+��E�S�%�x���G�?���%5��������(,pY�-�<�|�tD����7~�����T�&�����>*���a�%�}/� Jْ@��?aO?������U�,�mP���e<O|Y#��H��l���\|k�w���Գ�H�&��c� q��Ne��kv^仢�+�%j쟞o:���d�p"��w�A�"F�;����J  ��֢JH2����m �Dˑk����$s
�hJ����=�SSC���,�5z����ll˖ a��g��G���s�3փl�����''���+6�aT�JfC#�Ns	�:��Ws��?��4�.��g��ע��mQOE���9w�F`�9�|#����J�_�E�D�f�k��d��n�`�6���N�[���T/���@���.��^$�d��( n$.��y$yY�6̝u�Pi�2���Pi�M��[]���5�9�i��?0o�|_\��W﯑�N1�
��eS� RQ��֌x'�T�JJ��a�x���=`��8=�ՠ|�@7V�'�X]������71��;��b����!= Fw�n�^a���d ���8h	3�o"�I�=�����'>�	M��O~"i���Xs�5��!�)dyv.��]1��L�\oE��Q���n�]�0�����#�+�ƣye�>��OZ�;�}/�Љ71����YY ����[���t�9��f�� �:��!k���;ټ�~���D�|'��W_����FzffB�e�ە~�G<��7���?�aVV�$@Kf���4�=���nE�!J^��c�{���e/�&D��*$0p�A^�n~�;���w�kܤ_��r<��;�0��E�ѸS��V�d|��q�W��w�2��s\��A�Q�DG�)��@�T��:}�l-n$�3��$
�2-m*ٮ��ڑ����#�30(#Ru�mp~��3L��۟=eٔ	$�~��m�d�吱��0h��̗��ku[qzVM]\>��f�h�����uhs�ld����z�{�֖�cۇ�lղv�-��^��N���x67��n�B��?�����3��o|Ǻ;��0�]s`���i�~o�f�������]{��*�����-�k���x�Ϋ�����E�/%�}����_�a3���l��.�w�;݁�unW�ns���(c�DH8��g�9uq?�o���t6Åƹ�/�5�"Z"v6��ʹ��T"��W5:���0�j �7�i�=}�.=���CX���i�+�l�Qw�L��m�7(;���,���S��_<i3����ծ�`R*.�vy�G���Z�B{��ft_Ag74��[�s�ռX{��"�`�V��y�'8I�d�C`��ٳ��u����׷�[ϟ�6���KPB��.���7�A�T0���|"N��� ���� g�ƴ:�B������A�]�H���|���������09�3g�h?	�@t��	�� *8{��v@K0׏��cd=8�e�2;	�!t"� �3a�A�g?)�Ra���n�u�l,+6���<#2��Qcb<��kE�op@���e��h*����@1%�x7�Ը��$ �̫&?���Y߳�d� 2v���.��C�C�5�O���x��m�����J�"����E+E}��Dă\]	�>�ˡi	�~�$"ߍ�X�#����ҁx,������X;�3|UhPL�����lXm��O�Z�{Z�?)�(>7h�F@�Q�Q_r#j~7_1�|�( �e5���.�Jo�4*b�7d��S^ց"�!biYY�z%Hߤ��H��t�S,ː5�(�>=Y)Y������Y+�,�YVb���v7bp�脣R$�{D�Z,�a �P*���k	ٛzC?3D3*/������MKzR��8�@c �E ya�"n�b���C��*sj��:�He�A�5#�J$�&e�F�CB�0>~V�M�nݮ��O��F7�5���4E��ϝWetӨ���+�#?�����Jҟ��g��ܾC�#�<b�8h��b ��NTR� 8Y)&܌������5�r�nF�v�:<�ܳ�=b�8tH��jb���qʶ���LD�;������~[B'�p��`'��c70�{�ȑ�vʍX�&�+�@v��ƛ�ёazО��/UB ���m赞�.qCȞQV��*v��CD=~(��>�T}�A����=|4L�Y\�mc����W�Xv|��X�/����j�:���N��R�g�+���	0�q����q�t�R�ވ�
hʭ.U�C�
o/q��⹋�1��(�bã�� �!�
��U�ԥ�&r}-d7�G��F?[6^���+6qἽ���]s�����.i��>��(Q�HZ$L��$b';K�Q�h�{ؓm�"��)9<�A���;��?~�.�]m�)29�y�	?�p���؃;���E+�8HW�A���6��H\��&bx)�O�����rЌ<�R�j��ngO�c�~޺�l�3��y�u��'.��?��	�m��|���_���C u�US�<{9�]h4o.��q[֚w���H֨�Nvs 9oˉ�t_;�A͑wH�rú��|ك�3������~Z��\.��w��&�� 9w�~�� G��5�ٯ�پ��f=hs�Y��~t��Ҷ�Z��>��~�����JA�ï���j]՚6#Q��| �S�B9���FeMn�[����,�s��'ҶⶲQ�.I�<��9�kT�k�n���ܧl�� �����A�Bɟ��G�!�S4c��m��/@ rJI�.R"�3�M��}7qquY�y�W��a���^ͧ�ʔ���J�L�Ц~��e�RP��p& #1�3LS*ڼ_+}\��Z�X�T���G4�{��3��O�^��*e������LN����|��F6|��;*���u���M뺊Pr ���/F�/����q�62�Qt ѽ��^}��u�7l�g�ro��:8��s�t ?Uv^�S�7���?@�G?�q�eS����۳�<k?����<K���_��%���~?PHz�G2�}[��-l��x� P�s�ʋ�F�*U����}����m����k͵c�Ȣ�쩘��� :2���c966&[�ͥ�+��t�(nkoU�2��䓡��U&���E�u��0(�sgl	NK#%aWg��Ni�TF:����QR��ηc�Yyѧ�%�jR�"n��LPY!��9��<c�4	ڹ/�{Q�r?�_Z
U��q���6���	&�u������a,@<�/?��Όf=7C�]�L�	6||�Z�����A�oK�ۯ���Jg��xu-�xP4ue�N����J%�֤ҟx/,�hvg��qn8\V/[N�l7M���$%CFIS-2h�5��y%��ڈȝ��ux�(c}l��N9�x������&���	��?�~Y�T���36MVH��l�\[5.pU�Ż�:t�(7�@�Ev >@�4:�OG��<P���#�ِ��С hkK	Ī����w����sH���G?�Q-�:���#��K�!��g9rx0($�� ����5�g�Ʌ{�)m���o����։,U���`����"�?�'2T�f�8��ͰzR���9E�*�ґL��z����8�^���wA���/"7R���5��/7$��4�g��u:.h����}�݊ڞz�IeS)�mF�mR�^��1�iEFѣ���3t�ǁ��Л���H�=�a/��xb��G��(cJ���s��L:t3/-/){(cXo�w���u��-'���N�?[�3�Qc"3A 7֮�;�P���0��0���T�9��}����V��q_��m]�|M&�hm��V&��7�p4�nE����+������+��s�K��I["�cvs��Z�ckΝ���v[����Μ��Tuށf=~S��Y���Ҥ���������tڼ;�Ҳ��E
	��{�GkFSx��`��|�UTy	;��m�d�}-�6Y���>��K�߶o~�!���{����=ʤ�N���8��`h��૾��8�(�Ꭽ��mR)��R�hɹ-�����ϟy�~��׬ct��Q�p Z���
N��Qw�&.��a�ҵ0{\d�Dhj*����`�k��p�6�S!��i���,�������$�-��(!��g���f��hf�莴����P7{@�p��<�i�sS��E!��$�9��!�W��j`�����*k��HsI���:��_q����T�]�:��$�ğ�;p4��#��%g�Qg[�{����c�lp��Q 	A8g-�p&5V�VU�{$�u��y�9ʻ�@x���^X����N�5���?�
�_���d�p0w�{lˎ+�'~�L���&�$3��h `��#740QR��Fv�N���A(6�6�N����~�^��~pp�}�w��:_Cĭ�l�B�d���$]�
bS�p��nc�������4`�v��ۣ�cCnG�/M�����g��]�N=ol�+�f}Մџ��A�bU6 Of����_ػk��*�ؕ5������j~"����S*C!-� �B�`�Ct��0ӝ�+~�@ڵA2hx0����<U�J敨�C9\�h����b��5N����LDK(�ʎ/-]P����o���@!�'�u�L3�J^�&b�j�i�$�t�AP~�}#ԟV|��ZH֚��z�Xu��kFјH��ᭋ��T~1�Z�Q�Y��⹋Rg���\j�L��P�GM� �9P\H�!�O��]�H�L���f�����J$�	��5RDh��>)��#�ؔl&���^�Jc�f����<���h��P>-�3����*����k���ƴ<�f�G�"����VSI���a�I����5���l�qӘJ�_��הu��ş���U6c��J�qش~/W(	�]�^)?P�%�#�I$U��O<��9��@3(^��fAM dx7��m�&b���H���{�J ��Лo��ld>���mc�n�ɦ�މ�=�J �'��r=D�7�ڥ{�4Nf���o$���"�g�9��pTn���S���F�X��l1�A��J�	����X�"�&Nmp�O|��	 F�x~&��w�:otc�,g�}_A���?�.Z4����gR�����P�5͔�;�1$�]�O�]�j�e��l b�2Q=Ɵ��3'�gǀ#ѨE��n0%J���ڲ4=9֔ߟD�˟}kw�ي�`&r��N���c�l�5���i�`�t՚���*�s���jm^|d�#{��d�#�2�S��Фl���q+H:�==b�ؕ����_ئm��KS���O���q�2��9i&��Z��8>�LL�����]�Ī:��*C�L���z���;�e�@9����>h;��!�z|��~���3֎�g�ݟW��=0ȴZ����q�Y��� ��D��6$�]������ӧ$�m%}���������f�*��ElZ{�-��.B= �k���j����VJf�m���vlr^S_VȖ2��ڴ��`m�h=��t[�_+�O���h.c�`
6��
�%��EJ}�f�]'���.��n�e���<�����̷f���&��L�,���5��Α�GJ�`<8-�@"
l��8J�J��Ԃ*���8C�� ]�Q��GF��N�q:;=�l\&�V�#ǉM������qv��� ��A(Tap���0��UY��Ŏí_�j��*;eH��QnV&ٯw��=�@�
Nx%j��v���^~����7��M;��e�?�/L'q��`��ƻt$���[d�Xß=񄲨?��퉖'�o��ݷ�V��. �jDoa�)�� �M�g�&�:�J|?~�{$(�:�Õ���{���E )���\��ެ���M|S���;�!G2���slw�!��k8�>D/S����H�����R
"��ZP��K��g�M7�rc��Օ��n�z�l�}���I)[LMɢL{�zV{����qHz:{D-Y�@�w�~.���p5(e0鋵�g���"TLMb-�G�5�=�Dh�ߠ���g�΃�>RYvߏ�vv�^L+8��y���<I�%�y�Q�]��L��l4)&#u��dǓ+e��z�� Ot�i�W8l���O:&�Ъ�.n1�7�ƍ�t��f
�ఐx(J<���T31W���DP̯�/g*��k�5��%!���"�z��>�x��*B.�H6^2"݉����$2N� ���r$��q�D���v��ۢ'?��kA����:߸^q�.�U����t�ͷT������ѩ��ʝO����Kr� 	q&#�.;�,㫯�b��ۧ�H� �8�lT��2���G�y���l�nÆ�P�Lgd�Y'�(1 �aJgUZ�(�#��aM����/��b@��7�v��!�Kx��Og���32LD�n�)� ��8�A�{��m-Z�Z47�-*��b�4�`h�� �W�ܩ�UQ��]jD����uU�X����T�D� ��sMd�P)��f���uib�^���g#����e�#�Z�L�6��"XJ�"oF��to�8*:�F%��!�H�r|D��ާ�W*�rs�u��0�:��3Q�3�l�F���SqV}���i\e����l�����*��:UΠ�}-w�hRsF)�SH��=��g��_o��M����_Cɪ�w�=�14���!�/.XO{��}ú����v���7�ß���5��ʑ^����O����l�~&�7n�\�6�Х[��YBòR����8;e�5&��Dk�}�m�3��Sa��ª�ߝ��G>l�+t~��֏�n�6�Y���ڙ�i+�E�N3�����>f_����rE\�`�:|�5��_��h�U�N�N��3��O=i�`��n7]{�mں���kK�*�n�������)w��Nu��=t�ݨ8h�=p��6��f�9jCg2pgE%��v��k�ڝ;gi�ּJI�坩�Ց-����F�S�|��e)� �t��=���~f���ji���٠E��6��8֙�-�.=B��h�V}�h�J���t񼜹$t"�ed"0�lG2�v���R.�^בM��({���L����KT��2@0���*0��r�RDX���f�8�H��<6&)�.�H�PY����24g�M?�cE`oaa)҄M�o���K_����$����Ϩ�و�̀�����u�2[$�{w�y��:��5и��gx�/|SL�� �x4"׊*�1D��~�'¤�Ye�H����N=P�PM�����T	g�7ek�T����� $k�݊KƢ^E�����G�%����#���pU��1�<�X!"̈^��6ϛ,�o��o�ywww�6O�� ߈&h>צrrq��`Y����/h����m�k�?��xNS�u�}@����D�g�--_��A&(��|irB
�H([���C�psޕ���}�/�t?�/�AZZڢ�ր��^�~"���?De�S�Tt��A��z�>F�E�:5��=u;�L�U�5_������,/���[������Z*�e��I�J2��xeժn�n�a���:�,MY�o*�i}3"p�Q��`j�I�4�I����q����4�A�/V����XX��c�J��Vi%�=����e%x3����F���Hə��m�T�p02B�tq�8� S��t�2C~��j���&ڒ��jI�UZq�6�.���)�!�u�Q��Z g����?����x'&=r���n��{��㙧��>%b��>�-68د�C��gS��M��sO��d��d(����W)ejzB������S�9Y�pXS68�E�����A-�ub  �<#��x/�����t�Q� � �0`/����E">�1���|2�!Q����(j�+����y�l�뚚Ԛ�{����ݷ��jF<��;���Q��t-����04�3��܈��;��!��f��;ho�qH�wvȃ�G���r(�a<�>��Y5V�.S5�t��#���D9#K�h��U�М������VMeI
Ȧ������U
-�huR�d��R�(3��r�{|_��$s�UqSR��u�i0&�,ix8y�.D�[|/�-�l��O��vR��10�q@ZIZk�Uٳ�}�~����ؿ|�a;}�m��g�|fڶxT{�����v[pP� 2����u�s�J.ٝr99)0,���|��·L�bïםbr!gs3���W���tUƬ����G��]dJ��i�����_����d��d�6YY�[G����l��vfb����9��6��N�ԟS{����Gm*s��_�S���3hG'�l�xĖ�M�}�U�%j�����-��~������g�%����*�K\��'�g����{����[�C+��*ź�t�n��?��Ef���-Vm����_�s&T�%PO�Iv�	V�K*s���~i:�|{��������g������T'@������Қ~�Q
Mt�(Mu�����/4.K4�sj֓�_��6����)iJ\A��)-]��\q�`9ʪ�DAR�L|�t�D��v�s��L���^�g��>v�\`t	��Um`��2�kE���n?4Z�7�K@S�&�aܴa�$�%�4#Jz��$! �/���<:��GcŢS�6!�\3`��u�}����.D��Ujh�	*��G~`���o۞;����y�����ާ�y��98�_��������W����c�k���{�� F�"��!;����e�/ �	��\@����j�%0������}TtԴh&�ƙ6���Fm�ɋ!�^r[��6�kHEO�>����OB��A"�����>'i9�����)���#��X5���S�.AIۆ�N�,���V�[��Ԅ��6

6َ��ƃ
��5�m��R%��#p�V����+�݉�B�!���G2{1��ߝ-�&,F�2�!�m$���C��424 ���U�v2�W���B��" Y�����iC���}f�,�6ltm�^�ΫT������f���*N�Kw���f(5K��7�����"�����)e?L4�e�7j�jf`4|\��zB�S\)�M7 �/���DRQ��n9 �?�G��c�=�P*Q$��Z+��ͣ������������d�,��I��2D�I�s����0ٰd��<����9�ȓ�� b��Z=r��w���=�z��`Ǐ�����W�D�P�������� ��MnD،��[�0����k��R:���p��s`(A�t��[o�n$���_?��t��e�(�1��*(rya��|O�5���W�x/�!�`�w�:8 >�V�']l�o梱tDt �-�����)�G��H�#�wȋf"����Tc�o��E�<����}�A����tk�l&�Ed���61n�j�2 ��,	�?����Z����?��hm�(_S�g?c��;�����%dG���:���C9��L4<��n��/ȡ�'s��>��-E�E��d�9��[e�=`�g3jv?}�6�m��i:dA��d���{lF�����7du�� 
�����sn�E���4�ןŊ;�A6��w�f��%mmfź� �m��X�aay���f{��m��y�nsrm����
��j"-[��@C�\C�d%">5���H�-֞st�����]�d�p���m��g���BOmin�6o�M��v�܄�< �£n�i7���o{i����a��'�̕�(��R���Z���ư}r��ji��7a����~�����o+nm	L�>>�}<��,�u���������7��L��_�b��Hmxp�?������_~˚��@��I"���*:�̈́��@���Qn��z�,w�7*����� ����~p�P��w!���Q&����!��٧�&�\��׾.E���;�hN={���J��������Z"�� 9���?�3�`a��z���O2�\h�u'�'���Fp>8s�J��AuDz���2�-�l�Z���P�"��˕��c��F�/E���i�bc�dc7�) U2}d����q�����$�^#�t<ޔ
6�H�9�+�7�7�+؄X��%f�_�:�[F\?~}^� >��薱1�W�B�E����А�'�}��z�F��L��t|-�F�*� i����Qe�!`	w�k��A*k������s� (�B�/��e#�V*V�����v,R���咒�k�\��S�qh�::�^4� ��-g�;�����T1��I2�(�@A(:��gCfP��aTiL�`�Y[|6��ú�9M�����t"֌A!����q��1|�reeI|Y���+�0��+дBs(נ@�.^u�]�_U��Y���	��\��3�S��\Z6��@�]/��A45>� D�i���k2��Id����K�h�P��(���\-nZڍ^�RStG� D\��!�J'��6�W# ��CA�r8NN.��e(	�,���,BK^̋� L�	#��$�f������_{�?Ƞ����1w�,�AH�������6u>1�͉�5;)N�r�D��A�5K���������� ����Ҿ�_�������@�_��������?�AȹJS-��z��A]�� �H��3� d����[��m۲I�r0�ρ�N��B/�����Q��^' n�;��=�Ox\3e�l��6�@�b� �W��Pʦ�Ȭn&�@�?q�:�%u44�����{�FH��L�{1�}K�@g*���!x�0B� �q���-5� ��y� }�Ҵ��SA��I��߫.k��ޮ9I@":f8�T$�D��>��P����Ȗ����9騃7��bM1_t��K��HX�lJ�Z����U���9S��F��]�8�*m��)�6����8�3$��w�ixkA�FMX���|o/�/�ڭ���4��nX����O�~�3���'l��~�.Ϲ��`���nR]�BH���X	Z��N��H��헯�����G?�~n��F�Vs�S@!�٧�P��x�j��FU�
.-�J��k�_�r��4�T�5�=uƾ�-e�U���s��ƘNZ_�����[�l����ID��V�u^m�����&f����6�`mfy�6�^�����_s���}�t�j=��n~�?�iڇo�e	_�֬�ƪ�l����N�����_z�m���촂7����Nqq�P}Մ���,�񽞓�d�L���'_x�N�co�sk$[e+ՆQ4�d �u�iw�	��<[�	nG�iv�xp�m�v$f�i�t�ϫ�߰���k�Nq(�TP��fr�c=E6 >����J�r��žC�b$<F�f"@���O*A\;�X�1E�*P�n?���-�_����DRS����:*��>�|�^6;	�Š�& n��9�3�ߧj��m �jhB�r�gΆ*<9d`�;�3s�+|��j(7bk�f�����uA}J�P^���ω;x��i��X^;�{�Gu�u�~I��W��������odS	�iX���}	t*���^� A(�f�=�l!��]E���^P%�Je*k�t|u�) @���.~�Ѷ���;*4 ~*m\#B\Z�QN��[�>���҅��W�� x�<K�	I �@�o<�� �gnz��y�Ie�	ZW\y�:��l���kjMm����~���0/��D�ף�y1���Y�(�W�@�"s�G2�q�8�5�Z�X'iĠGAw��/ ������I�+Β�EIt#Ъ�ϵ(���c}�V��e��k�L����*{x��(ۙUN�	��{��h�l�L�ˌ��Ђ�/|$=r	Y�&P$v+0�.�P]��2a}�Y�N��]���RU=JfbC��0���O�y�LNY^�,�Ē�q02����#uu�D]s�� �YŐQ����'��5����U�s �? ʏ�]}z ��A�D���i�Q'���?���3;;����7�@�&R�����?x�t��*j$a3БG��D$ݶd��D�\�)����=������X ���WD��ۿ�<���]wޥud��=�L���E4��ᾈgf�Խ�� w߾��B�� H4�Q|)��3sxO�:�>s���?w�~��*��h*�����8�?��f,tN��{� l�e�������{��3L����'8�Cn���X��ƀ�o)7�<S ��֟��n��?�ڟ���n �\/p�j���>����� Ŕ:x�Gx/Ȋ�'cLWB�"�iMpD���uE�l)�t,�N �^ƀbD4��ח�%|��әt&�fִ� ڱ3�s*�I�)_�r��˧:R�g݉����Nڕ�t%ǵ�lٖvz.�5��� M!��AѪd��n]*�m�A$z�]n4An���&�,-���a��Z�������߆�:�J�>�����W��DGp��\7B�!j_�����?m������o�����%�p�I99������d/��2�	���9��|E�-�&�x�ZZYS0y��	�z�;���e��wHy(�{��4�J� 5������+^���V�=�ZZUG�<�M~}m]ݶ�h�T��;$;�sӠ�OV&�N����C�x��pk�!3Df���<�����YˎN�y��-Y��������ղ��B������>�M*�i/��M���Y-��C�!�"�;��%d���Y\M��M6�����o���\�}��
����di�|��#�U�Ɏy�a�&4���ѠHty �)��;RH��sy�P�R��z���c��z=tT�$t� �8�"�S�m��S���`^g�m�Tj*��%���u�������a'Euʆ&=�;�SՆ�neq�9m��i$���b�y���I;�([��O� G֎jI�(�J�F�K�b� �k�?���~��DE*!TEp�p�ŝ����_��%N���]�u��;�D\3ώ�! p�v��ݷ��n�5�M0�D�o������̮���O����@l�ɐ�?�� CQ��3��3|��j�!���� ��P����w��C8N?a7�r�x� 3�E���o�o��E	*p�Li������ �uN<�V�7���^w�yV���k���v��y�Bv�&�Ip� ��T-Ȕ��Alw��G}�F���U�գ�kZ�ƺ�A"�o�nq%#N=��������no,Z�u%�,C�5���ϵ�!�45�mW��V_��G�P�zP��xcR����%�Z)4�P�M��LK�Zp8;6�Q�J��fݘ��`����Z_��u�5�~��K)�4B
;�!6"%~�W��Mtɺ�w�s&j����������D���$M�y}��G�DA���=��!�z�����,��&��;���l�v�2��8�+24i�D;4���b�`�m��*� ���]����?]B���O�{�t��87#���D��W����/�E�-����f�kn@�C�� ����ȬW"D�*�#KG����PW���2Fu��^y�;��	kq@�!��>��GZU}6��ﻱ#��hk�M7�0��0b#7�=�݊���ۢ��N�e���.y�5-M��.۾#��ۭ��d�>���_r�����A(%D��|��{��^�g�>����	(�P�' !�'�A��}�,B%Sq �&A噙�PB���a�)�ʹ:�-��Ô�X?������J��� ^�}���M�Y������ ���iܤ�3 5�I�[�.�p+�A�9�V����G!n��ɉIeK��Z)j���ʙ�|F�(6��hfi���+��`��5,�����K�� x�	*~���.�Y���9$	{k|���+��{�,��b�L��s�څq;��o�>�	�n��/������4�h����]��W��}r���;�5���q��Lω�lu�~w�͊�茟��Uܨ��ng2mV��J�U�F�T��p����P���������~�h�V�yM-�Z�T�|����_�C��FZ�ōxZ���������a���,�+o�>��M����ɺ�:�ę<3�lc��V=1~V�S)%���p=��4�4�����V+��|�m�2j�<�<��lU?W�|��6 ����?n�z�n�骝j�I��#�[Yu'�4���Ξ���]�[��?�����IK�ޜ�=��祖��\*@ �fDH�=Ld9୻���3��Y�]7l�E�Yː�]?�	:˗���UM<e??�t�#���`sɢC[�_}�̸4���=D���x65�s��Eӎ�j�ȄLa=J��5l�U�*F2]�҄h/+��s�F�����_��J<��s  #��a;��J�2��(�_��J�>q⸲X�l�wŅ��`��<������H���D�-nk2K+�-��-|��-�4H��&hNy�!��Oʾ�����;j� 5u���p����7$y����4j��'��}�fû���9����k<p�*�����)�1�Ex}4�`�HF�q$�	��~%�����4h���g4*��PI���1y��)e&y�e2����ȿ�/���[(����Dϟ$eydx�.��?{F�@9�m�o�qP{����?��iqiA�*8�7���5������V��l	���6�8e^�W��R����v���:��@_go��رM��҅	�����G𿇬���O��jj�a�ʢBmXo(�����ѐ�/�}cA�ta�]F�/�??f�'�ِ�HՕ�l����Y}%ɚ*����i��EŰ�#� ���L:� �R|�}O�B�+M9,Mc��E���S�9���6�p���#��v� A��d�:܁�סу٨D��sØ��2j8D�t��͠�xoy-J5*'V#�-�f�Q�`{:��3F�I�52�|FT�t84q�
������;vz�uX0�^J�C��X����.�8��d(� �T����ċ1��Ct��Q]_\r][Y��+������ՠ���^Q�<S@�9�T$�$K�ADf��Ɂ�ˣA2Zd�(�8p@Y�x@��5 ��{G��kJD�7��sh�g�����K�aێ�w�:�O>������!Y->`�	��ƽY
c>$������(�H�����������%�-�@�32���5z���.G�>��ɧ�T�zϞ;�ـY�&�ʒ=��t�Uec����� ���� ZM �mѴ��iO&X����pl�(���'��Q���d5prp�C��k'�L���b08wdÔ�Z$�Ժ.��a��µB�HEB��&�M�>u���&���b�b��F�`n�r�wW&�7��Ux�=��~������D�¨��ظ��^+-/��?��=��_�P]���|��-VJjP��9������~�c��7n�mL�!|���*��>t��G�c�����ܰV�֝n�	�&�Xe+�Z-�,�����\����m](u��O�頪ſ3��O�8P�K�"�F����5��j�����I���ђv ��j�J�	g۟˄�Ţ]�@�mp���`�E���`��W^�_����VW}�����V�,R���L���-���Q;r̝Ck֖�n�{��>Mf!�bk\���/~�+�{���[s��Tv�uؖ͛lae�f�y,�}M,-[�׋�\u'0����LF<�H}3�E �n��⾗_s�d�ڑk��[ɟ�Ȧm�<?:�ݱ��l��p�ø���,T��)˃����0})*�g9��vb�����ﱿc��l�ۣ��NuvB��5׫ue��
��� �J��Z�Q�O�x�|w���3g[<`�3e��#�x��/N|,/i���Sz�L���WM���{R��q�Gg����_jl���w�]{�u*1�V������|��n�$����1v��q���{�N���\{M��k4#�� \��d�s���|���G���O( ��W�bRi�O�D����X��Jԍ7ݨ$ ��.��\4ţ�ם���w8��<\�$������5j��'��E����_�i�&4,ak��H���?ɐ��Wt���^b��(B���j66�I����Jі���/��,��u���1��I6S�����ϸG�r84(�NO��o��v�=� �g����k�^T>��B�.,������(��D7��P<�0--�{��Ɲ�	�fD)�\���GU֮�u���Hr
H6���3(,$�{_ӳ��hV�8W����0"�M����_\̅��l�����,|@.��-�G%"�ZCz�Ef��5��:8���B�U`0B�&�,W�D*#���Z�
w���f�����2����D2��#AI�� vww�mۺMCW*�i1DNt�JnG%�x �8o�X8�l\�C�(�����������O}�r�߼r�%U�d�G{T�����ܾ���k�ߴ�|��yċ#�}���/Iچ2����޲E�����xt4���Ai�m���(��[��m<��ݷ��?<�Ѿ��?�g��Cڟ0�P��ﵪ�7�	G���5��r�{���W�(��1D4���䅨�B��T8�p�R�X#�&�xJܔo�R"����{�[�
#1<<d���gu?{�gfݝ*�PĒ3al`s}�F#�!Ɛ�6d2�"���\�.9"��\S2r@4�������"���ᓰ ������#��� �x?�ZK��y�Ȭ �LrDʧ� (�a��0�W�2����hɜ�\�#�l��HI lt;rܞ $��%+��d,O�H TP�ĩ�i�~v/q���w�JY��n�fM��D�%�j3+��:���<�Z�M��M{�V���F���&��&d�
�~�xך� ��-9(m��V�>��m��Z��*kS���XA������K�����\d&��{#�siv��KD���p�F6���;5�k�j����vX��1�)W0K�R�dO�b��k&�h�#3�7���C��T�'�	��,�E�K��������T�5�Qz��S�sZ{*0%�(u�33v��i]�8��3��w#5I�I-R�X�s�<G�hGb�HcdyV���t��|넽}�tq���p�6���֍��M��Go$�����* �����<�A���!�h�.-�g�)3�/6C�������&���J�jJrQ ����Ʒ�E���
EL7��=�K+Y@�4��lI�*�M��ZWO�ʗc��dW(�ҹ��R֧����*�
�� ��- �a�{>t�ۖ�v�}�k�6��N�v�8qQeT^p�n����~zЉ(	&�	�iRAu��{u�=۸܎]��i$��.�0��'>�	����t����~�a�
�XY���Q�i�H��.m�PyN�	cNIH�/�Z(���*i��yG~~��X�ɠK�C�.��V�nn��}�Z�\��MC#	��KTeA��h��No�mf,��gM���⪝��P�n�`W�R��5?uZ@���f�!�?\�EM#���Ο����-v��9U����L�#ғt�GXC�)�lj`�ng2�j,���9)�]��)��0P#$��|���������w��U4�Q��3�������Hj�mO�2C��xo��ۻ��;���Z�WkF3w)�cr|�G�	źdDv�M9��yI���n��:�8p��Z�к]�n�a�/�騃Yݯp�[�F�! M��ډ�Hݼ��aF�:64���,O���r���R�,4�#d�D������-�@^� ��"ey�$-�`��C?�yL�]᠐�*����?��*+��o~[I@F��w���Jˋ!��k�ӟ>�C������w�^�/~����Jw���q`����P��D���&�5���W�p�2��Tv����hC��x�]w*󕌦�`�0*>�pO�'#�Mi$V�G�u2:��� ���$�zЍQ0�	�k:� f��a�=#�$�ea ټ�$�r�0����2�d1\��P��`�i�ãRx�<C���{b?��IEi�S��e��9K���$�̋F'�+ύk@�'��[<�н� �����BdI	:�RlFN:��� 6�QɈs��1���gb� �0	�74�<�|^5����3�hQc7�G�."�3r�����V/��y6�$�4�N���5�N2&��k�;�}�"a�w�oEnʅ�b�J��pSc�V*������Z�;�fm�Y?��G���ΡK̃/���]����s_�<�J�iݐ���ЕM����3�a�$Pe���lZ]ʭ��d'�� ߕ��k�M)��E):�bh@&�fk��j���������i�u�iu�p$�����D�I��%�u����04n :	 r-:c���R�,��{��x�:��/؉��\��>W�~<Xmb+��iJ�{������ I�߷��j��w'Y�쵕x�M�����ݺ�*�:?n�+�U�
�d��j��y�"��z4�jR�E��hS���� ����*VӢ����W ���Z"jf� qm��1F~IM�Ȅ9�ͨjC�M�ݽ�4�റ���ќv�u�Z�����A/�F ��;��t!4Нu ���,_�{L���|E���K���1l�6�e�n��5$:�α�%��&������(�(�|,k� ,x�d�����k hb+�rR1�G��/�;Q��A L��/��c�m۪���H[�%���TxH=���/q��wu�{���3}F3Ҩ7PA!�&�i�)��1�ŉ�c���r�H�:�k�������\c\�vl���e�bSL5�H�
BeFe4�>O�����<3�%+�?�1�y~���������V�$���)���=adL����Fv�ǀ-6���w�!�]R�]U (C�kU��}�O�O�_L��l�������c�y'��1�9��b|��ׄE��,ͿI�/��w��y�綟�E/
�b t|�d��C��į�Sa��\�G�t� 묮n�ѱa2M��������(36uC��OZ����Qk��)�NfPk�$e��% ��A��,Ϧ��1K��{Ns���Q|.a��w��{�H��a)T�mc��&��� �i��S���#�K�."+ �Lڪ�+U���T!֎N�JP ��ے�����dwg�P���5�I�ˀ�]b:x z��M���"� �����I�.Y`��q���ĄWY�)��0�+��'�EG
3,x��!�U(���B(�0/P��$��EQ�f� �*�h�\ڄ�&!O�;*���ͷܢ�%�\��(c��S�?n��Ay)���)�d�\x���_���%�bܶ�-ɰ4�y��<NQR:FO�a��W^Ea|<2�:�ʗ�B�%�0!�y�fy��������������"��ħ�t� �� c
`�%N��ƅ�^(|B�֝�.\t�E���*�At���T_N"�HE\z饑�iW�-���.�?a���X�0�Dt�lTеy���n:Y�4,T���������^�os��W[���"7��(ZV�)�[20��A�OM�cʛ�0u�I���⪻K����I�}N�w`1��7<js��_�a%WcFhJ�Ǭ(quIyJ�ќ5{6"��;E�`n{X��Z;7�ᩌ��l(Si2�*V*vD�&�y�(2&���H�.I�&��Z-���҅D��(Y�h��CFk�����Īd�d�������I�U>��M��V��a��p�6۹6�<k��Ł��б�(c)���jA�%��&������`6���1���_� �KS�C=��J*��;CC�x���e�Ή�D��e���p��X�XYY��ސw�`gM��UR�dpl�D�ㅃ!v�BR�2)������d�)A���^�g�c��0*T��E~�4s�0����})�F��<-��TcH������B6~М�V"gpm��&��B�7Sw����,U�E���Z�Vū���IT�9�m�lF)�RյH{
1� Y�)��'��q���ۻJ��A9�%,�ٚ����*��Ez��jYQ����]:(���Ut���Vxw��)��K�57�{�ҡ,�B�ݲ�I��iA [F�@P`����m���(�7vX��λ��7�T��5��rꓣ�=���LĂ4 ,���T��n�Z������c����c"β� ��̦,0�|�}�@
�N�E	~��|Lec{_��{a��N�[s�9����i/��NX�V�]S�t��aK��)v:�>�	J�߻c]׳Cy"�H��lsd�= >��cJ�b[�����n	'����c��d� R*�2��VhU]6�=�R��́����o ���j�w��S(b}sg����*�a�>g��Ѭ��V�2�#j�h����<V�έ�[�B���Pk*9��߽G�r�q'h_%U��-0;m.)�%�����wx�Vs����%��\�'��}(��gT#�n{�?t��ٳ��9�]���)8��P����|�?>��ZH"[I�����c� ]E��-
p��5¢�(Ԉ�cap��(�����ӡ�j��&��JL9�E�O��Y+�[ĩ`¼6Y�r( &g_��0п�@���琍���D��5�K16�PR�sxe,\�����J��� ^<�h���~�M����3^,�e������������\n��E�}��i���Z]���"��H�*Ƽ*
 �{��\1�/��2	]�fc�}���hB�������\?q�*������K>Rz�6�㎱!@#�JqUۯ��	O�O�{a�<fe\p6/����.׎"��{�df7�/���U�ʐ���d�%Ɠ6p�OƆw���)��V�,����I�`$>��O����b�<�~�iy����7)Ƅ�z�,'���DNw��Ԗ�{GDve���@�%� ��73�ۿ���)���!W���<h|�2.��L.v���7W�������� ��.\nבh��t�ܙG� �J�#�P�76�B�$��;4�������+.��0�B�eF(�J4'V��jq���x$H�Ӗ�����A�E�#�����x��2\��V,�ׅ�O4��m*T�S$Tҧ]Z&�4ʨ�@�6*�)g��=d���O%�K��10OeS�X��s)���� ������AS-מt��K�4*�U����l�pRO-��L~��4����2`��B&�Y��=�"]C���hG�X��>&YA^�w@F�~oV�S�hDh�A��ׯ�}��zG1%��]���yI)U�=��6�� ��m,U��|>�CcP�?I���#�ŹI�mJ�5��-ը���D鐔�*4���
ۇ�y{�v������EW(D�t[�lެ�(�F�R�)u������N����h�g���7����ʆ��L*/���9z�&7`p9��΅$����#G{�}���=������ʖ��x�2��#ڻ�M����Ml8s��ie(DW��Vp`S���"X��!g|x�#n��0Fn����}�~ݟ�sN; ҈��ɡ�*�J�hB � '�����*��}��QԽ��[x��A���u'��}���7��=�'��E���K�a	��|�J�v��=|�� ��K���1���?��+��!�H��*���ؾ�ŅXzW��Uݻo�W��=���{[�d$Fu�d3��dM�������쩢E�]Z�p�:!/�B�fr��E����!i�j>���S�i,��բ|�z@+�YQV�Z]�l6w8X5��9�ȇ_p$Ɇc�EYp�h6j1��}���ZE-��T��s&ƜEt�r�������e����h
�,�78'鴸A��Z^���H 9O����U'�ս����'i/"oь����eしE��B�s�R�b2	�ۛ�]#�(����d��5���O�Gl�ç���K��C#�#����A<4�b,`>�+��B��F+(פ�[slx��GT,s�g@2��o���'�"��7\�z�1L�s��a�c<Q�W#v�:)�!��22�D�&x�͛i�QS#s�=k������8�˗-�{��)<�}�C�w�� >��	E0�����{o�F���o\�/�������y.�h:�J0UTWc4S�R�*���C5 ��x0W��lk��1|F ��ƻ ���H0D�X����$Kdϙ9#M�V�tL�~g�9w��H�95�8�)��)2Ro*�2՘�hnHOq�ǭ�θ�P̄�cS^
^�_��g�j=h&��H�D�H���fUQAa6��\O5m��0`�(��g���0X��9�}!?UA�Mp�聍��܉�e�@N��Հ�XL�����R���{TW bZ�yOլ9�u�^�oY��CC� ���J���Tj�f#HX�Ǫ�G���φ�Ni��gc�1i	ηt�K�Ԭ!�|B���r�w�sx<��^�:�
4�2E1�$��~D[��ؿ�v�1���1],h�F��2~P\شp���M��?�`>���"Eo+��b�|(Ǫ6��4.�c�k
>`-��e}q!��������4$�l�dX?�Rk5 ?�u�,��)0�dxۻ���9=}r�X��gY�G�
G��$~�ُ7�l�= ,���FP�n��_|A�_�(߁��F*6�,�����si4�q��FBڙb���`����M�ַ���0�)�sM'/������2&����<r١R1��bu��wt�sN/^9`v�-Ej��M����^9Y(h5��{f����pOw����Qq��D5�>|�=A��t}D�v�]�,Z�����8�{�
�=���+�7�f_�5/��=��
�R��B��06<��;˖,1G|A����.1 l�~��0U�r�K��Ҋ�~=����&Ћm'e��{�9U�>'pd��)J}�yw����1[�۶mo���)hѾ�M�7����w����T�D���&�l����{&�\�YsM����Z&�l���%����嚽|ZD�LN�T�I�1kRfO��0wNo���L[�!�q�%p�� �D�'�16����T)W*�?K���Pr=zD���vyDB��+XA⹐k��]�v+��F�}A��vT��(j��V�\��5���r�i7J����Er^��Y�M�,]��%C�v,N9���l�W�`l��3��\�a��7��mM,�؀,�ܺf�	�Ҕ@�"�P��.��"ZƘ�qƙ���0O����/~1{̚��]��d$vR�$�}V;�	�d���	 �{�YMN�րDƖ.]"��"]OJ�Kj��7}SƋs�.��ɃF������ m��w��BOW��^�zs�{y�/�-�e�x�-6P��᳼/�H�f�XH�T���x�*zf;`.�G?�QIT`�X�ln|7�S��Uc&"ɜ`͆��#���[47�$�D�����p�� &MO8��cҜ��O��0�� s�sO��"�m�����Pf�3�,f��_"A�fl�!�ȅ$J�ᙄ��{p"d�rvB�ÛګE�R�@ϣ�Y�97��Z�9�Ji��ـueL�h����& ��]ebDM�O�6�LWEܻ��
�U� *����S.;Ϳ\�=�'!ڜ�U�W�	��0�Q5Ww �;42��#`��f-�E=���/�6���)#_�h�9���g@�2F�����a��!��O�����k��% X���9��¡�,xMm���Q�E��_E(+���D�(J���F�Cg�.������u�0Kw3��5���W�w�A���5����ȚT5<���ޕ��k��U��@ºa=QT�l�{�ZF^M{F����6�H]�H����(�O��8�k���r�N��KLUTDA:�ds>c�c3H��N&j�x⤲��<�,/���L3��Q����zw�߅��_�E���ܫ��9�B�� ���Z�昰:/�U�_"�d�H�8�6�� �⹱�lڔqj�V�K�]$�^�f'9{$Cl=����bW�"�g�=�?3.D��7��AY�p��[�|� njǛx����Vl7��H.v�����rR�����x���k�q�,��7��=�|5y�ԺR��R6���
����9��j,��;��J?w��v�?�A:�����r�DZ�H���ʠ����C����36#�E�'�|'u�I5T��-�2{�������@T�����d��&�&�}��P���!v�s�м$���A��M�9��(_�=h<��bK�vR�`)d���6)�����js��-��f����	q����f�tޡ�A��ʚ�)JT� B}2LT�m�R�X�&��tn���`�"o��Ke����2�i���C�3��K�̛'���^U�%�Mbwxy�l�a����S����!�V:	mba ��,z^*U\�xI^ii�9��g��A�29Zb��6����օ����c�&�-?���<� ���d9`��M���&RD��#/�C�Z`���C?'�̳��-н�A�~� \�����C��˯�\}Mx��G>~�����=e��Ü��̻['��Ș�b���<8(�A}Am0).�(��D�޳��s��,��Ҍ-��c�7/�$��C�{vo���Hd�S/�Q�n6�sSp���`��-x\|Ο�"��ɫ�H���� f\�B�V��X�3����#@@�t�ND��ف?N7����DT��K�J,by��<E�XR�:9t���om��*B��&oч09�/�u)�B�%���l�BRԉ�x��$��r���.#Ue���C^AL��{w���� Η�E�)����%u�r�2R��F��ek�#���+JRւ�Q!)/?���#�L���1#
���t<t�-�T���1�G��H��X�����0�jըA]�)�+V��	q��C&�4\������5g�$V�UB��W���9��p�Jd�ʧ�g%夘j�)>�޵�1���k"z�f"�cV0�N��	��JC���<���"�S��ڻm����a��g�6x�S��[U�Hrٸ�9��M���uy��#a��D˜.��b{�63�")�"B����"�*la����9�~���ٽ��n/6�|	���#+{�$��Q�L��i���V�(+ �$��_`6	�}�F�7�SR�
{����5�U�Gе'V8���^p��HyJ�1"&/���1��=zO�-jJ�����^������s�JT�G��?�S٣s�=/\q�*ȃ�Bu2QBh2�e�9���Sj6f�z���4�D�ٜ����a�n�����ЖM,`�b���}���Wu�Qa�9ؤ��`��)�@��h6�O�f쯌'�w��g����3�מ�.�`��
m�.�p���bk1\t�ELD�&�y����M�dW��"3GT���}�5v���1�S��|�<�ށ=���d�&J��,]�P�����P���h�A{G.jhk���C�9x��5���͑O-#�(�W�l2�M㭶εw�H�
��30����(�W����)m��!�e,c���Jlf�G2lj"�zw�z���rA�F1���E�u=0B�kO)M4��P���j���BV��K)�o��d0YX(��2���e#��0!ݠ"��Q��S���AX�U]�7dfx���2yZY���@\{H܎)�8D��#e��CQ*A�]1��Bی��5��W*z719&��LZ��C�Px�pO2�L�	)m�mL�lW^��=j�>���N5:�����\F�|Y�LL����/��a� o�Ϯ�A;7�_ ����0�o��"��/���!`���=����8�_�XƖ��$�?�}H��q<������'c˸�?��3�'?�iXs̚�?���(>0���-���7d�0� b"����]��w�ȸHᤴ��.�Hcu�����n�n�k��}�^���?���"��'QQ1�>$��$3 (�CX�� ]�KI@��$ ���_��=�\�gN��j��.��pb�0����b�1h�<G�U:�) ʘ�ǉ��a>�3�mj�Xsn-ix�m����]T؅S��g���bD�KP�.��J=�[}!��H��\�����27˅vŇT����鵕�<��)c�Z���P�Ւ�b��\���6�f)֕@�4u"v�DNX�n66{��Y�0Ʌj���k^��y3��*\=�]��6�w�e��c[�L�Df=�"<�_U$B$�+��Q��  �ઘi��pU��QId;Ju�)�� `=�MkQ'=_V�J�f��ě��x�����l��N�� �qKWTUb��*b�q;�}V�2j��c�/L�Ec����4��N�h.#�imM�g���r�)L��H1U��56��)��<�U�V�6���k�&i�(���1�e����O��[��9����S�3�b7ޝ��(�
�4�k���
]�oNU��اu8�۳\�q"zc�2��ȳ�3�T�"�����rb�c��*Q�׭���� �q;���97�r�%�� & �%#K��jC���{8�\zI8���s�;WT��}�k��D���6�[*&X��l F���,��HٜǞ���S2>d;ڣL�]]=zF�����9�Y�N�={�M��r瞪c�o�)�&Ł��~ ���r�@;{!�S�F©��W�Qak�=�5~�^y�䓟�}eи�s�y��·��m��f<�%7��
j�W��j��L�=��v��<�=���I.��;���ֈ��I/�1{���Q�7�����7^ؾc���]��7ŲR�15�6�;���R"���S�;�^D�@��#�mϬ�B�l�C+O;F1cZ�{�NϘ�dS�C�w�)��0�K�G�)��������xd^ב�7�=
`���t�mQ��}5sB�"��[�"���oK�Ir!�b-HD�i/"(N��Ƴ$� �15,3[�Do[a�l��n>������P�6c'��|�r�N�����I�p� �{u�"�����J���\��Z�JC��c!���D�e�"�D�H%v�Vm�E�}i�{.��b�����+>�]wީ�ą^���
E����E���n�H��D��!�Z y�T�Op��O9Y����zX�A���v[�D.\�Jh
��3zrq���a�Z���"%������!�G���;��k	c��>�~�uMp��2���Ѹcケ�f��8aTN=�Em�ƀ��K�b�� ��{��F��jU�Bq	"��X�t�O�S����� 7s�#X-D+�w'-J޳ҵ��޽��(��R܌���%�$f ����Bj�����$�91�*�ה�cT������cy�c�����%��5���]FI�aHm���i�e����g$rp�Z^�����f�����i��<8��:��E�W��.�_�0/�x7����#�^X���˛3Z9�5S�`R�;X̤�o��T�&=�p��E��a�TO�QL�nG��!�����|&�p3�Rd1�x�vӸ�#�i��Z�5�1�m@�hsa�@�����F'�����v;okW�"��;
x�l@q3@Um�s�d�'���҅��v�@�(���Uo���6�0�+�H��=k��E�i����6����*SR��]"4�!����c:��TSlQ�3W�.��\*i�TdR]�Z�'�.%�S�zЌ��L��SR��'�f�l���h��
�́޺m�6w��l�VR���M$o2vOQ�)�HZ[ԁ��_ ��{�����b] ���-��7^]�a8�W_��JT�����o_u����_��;�A��e+(y���4��]�W����Y6���<#\������x]��D�%l(����y׮=1�X�"��Jz����DG=�����g$;�����&���~���kh�r�d�2�)�*0G���) �ϓ����c+K ���c��Wawi���ۉǯS���2�N:�P����;O��&����gm_-��D�k��)z���{q��6k��� BȞG�1�w���9���`��슲y�(	��������fB���E��*��g���z:�Ek@�vY6�(�А�9�.�~	'	+Uc[�h���	����6��$~;��@�|Ԭ��B��Z]���*��M톆m��?�T�*e�5�D�+�j�L��PP��5	C����
���{fU���\���������<6r�s�C����J�>#G��Hd��{"�
�.5��I^��s\?U�R�����vN���РU*@"��ؒM�z�bo���:+��@����0��
{����K��q��}�c��<��\�#�|�-�f<0xL�1<����4���YѻSO=U^�JtO<q�
4��?y�'�e�ȟzC&�ԣ^<C� ["FCt&��z�r\q����X�Kl�_w�߅�_yU�(�ra����%
@g���O�S�$�~��н �������!Q��X�!����駟�`-cХ����!���uk%���#�~β{����~X�[�Pyz��,bޭ��6K'?��4��D�G� ���yRh��o[�`��b�������/6���x/l8"�S=�~J�QX¼S�A�N�ٱT]5P�����hq��h�I��We���<I�FǤw;�2	��@&��(�?�H�'"��N�NM<Cnn�ԵD��[cyЫ�y�Ck�ԧ��2�2�������2�1�\��<+�|U�H|�������f7�sG߻/����TQ�fx�H9��р��( 
+�0���d�Q�a󳫥.�*�rA��0#N?�;�x�G��*b���d9̧���5��#DK��/ue9(�7��'R;�EZ^��z7l��{�k"#P�W������M��Z����`ϛ?/�Dx�(veJ�p�^��N+1� ���k����qn�a��Y��7��gc|Iú��F�h 6�(!`���Ud�޶=��g��ZF��E��]�@ ����, 4� š&�ﾽy���w y�o���+|�=�+�Gm�X/d�ǉJbkj�
�P��[{�A�<������SN>E*!�I�#b������b9��r�hDDt�l���������5��x���9r�ٯ�j�J���
�=����7���������4i�d ���;0���*��`���Ȧ.q��Ǔ��rlH'c3ٟv��\���nutv{`)�m��XT�����W� $� ��K�hH�+�����w�)|�+Z�x?�G"k���Z-:�`�k{�͕�>34t0�u�J��u���D��u��l4p�3��ev��wج"���T�x��>�uI5�Ǖ,�:*�Ӕ���B�yR
�����4�C��<y�x��C���1%bowhio�e�-��45��*�Q��yo[c����]���s#���l�+�fi�V*�ZHDG�Pd�/Y�L�E��'���D�J�~k�ׂ�� �?��O4�s _�⋛��_�=�xE� 3_ecO�\��Ԧ�{�{A
���^V����Dʸ6�b���mb������s���s��ߞ����>���s�y�x��Q�X�O>���r�m�` � 6U�ޭ��Cq̱��� ]�mL��a�p�m�z�;�>^v�e"[���Q�B�<;�<]ײֽ����o@&ա���+F�4��q�B�S�&�F���ㅒ���1�j�J�X6�O|�����ѧ6W��J� �φ���~�y��zGD�|�5O��8���\���1�S�:�t:�s�Im.�wW�5�Uʺ��w�R�*w���N`��9iރ��{D����q�<E=˺���I��;�"y�h�L�~��)`�g�3�pF¶�Xi�Ii���:�;(L��(ߑ�S�9 �Gٕ����,WLj+Д�����i:��3�;�~cc��Ãn~�����EPT1�"�<���Td���Y��1Ǹ:��%)gvS>uI�0����2z�G:2�2~���r���8j>qo��Th+6�=;��<lN�j��c|R�p�m�3o�8��ѩ��8lʹ����<t�g]~IX���뤖�)5����({Na�9=��@�E:�T4�0���%��^��H֧�	���>��w=NtwSKK�Y�sl�����H�c &i���E�尕%��-\s��H�7Zr�1�6��)�ٲ��v����R�.[".sѾ���6~���9�-��)��t)3�YcO>�P�Ŝxx�|>#�L�@�m@�|����8anS�L�� ɕW])���CT��p�G/[.�X�9zq�jr� BD�_�ֶֹ7A1��>n�E�Oفt,�6ƕ~��Ұ��W�~ZϲF�(�#K��2��p�� �k�\&�|ՕWi{�l*�V�Cb�1`s�駅�Ǭ˗���|��d� ��|��Қ�c���k����)sHe3�^�1@}�(��غk�x���Ǯ:6����4��iK�\���DњT��.�D�&(j�w��{xhD{2�H�c[Sʙ�rI��t�S�33E�G�|m}s���-ʅ:#N���/;����������gs�\�_�߱? ұi��?yJ���*�mޒ�TC�]#C�(}���c�D�i�%�B� Rw�R�����c�6/��]F	.ul��� �Wl.ze��)W���7Kq|D�f]��I����'�����p�Ѧ0+�x��:���$���
�t���xʱa!�y޷����j��<K��e�]�׮�h�	�=��*�Q�SF"���m �p0It����pO�B2���Z�<Q�o|�p�Wo�v<��~����g�\��ȸ<@�2\E�z���T�~�7	�^��۶��Jh"{x����c ��w� 5i�&#��O:Y�ṸO���?f@�l��c�X���Rᛪ���A�8F�����[����/�(\}�52��\�˗�E�N�" Ȍ9�Cܷ�<E�z�*�,� bLy��\�χ�G�������O}Z���iT��˗/�_�h�{�}�]�xy��E$��Y��������S�����d�!���46�EQ`�{�7�0o�G�g����a}�Bm�����<ډ�����N�p�:�����.��`�g��%`ځ�[��E�%� ��4�tr]�8�#4�Q{_c�v��������[��tx�󘩠 ��a�T��̆N�Y�L��d(�$�%ۓs�'��a+J���%oTP|ǵ�3���:S�L|@�� �"2�n�I����jY��&sܺ�恆C��f6rNWG8a���9s��ѹ��n�&���BWGk��&�� �9�h�"͠N�����a�A����W��j�v.X0OŌ���L4�J%Fx#7�he��� �Y�UeP
զǘl@ol�k����p�������b#�L,\�+�~A�9���Ҽ�=[ɦI�	E��fϚ��n7߳����/Gڏ8g�}���.���3��	���k�_w�?�V��B�x���$�q� ���lόM���Pc��2���}� ZH��x�7�.�^�Y�{��R�hn�; �8s�b<q��6�9���S%��?,pˁ�� ���F@��NM���DS3FDAm>O ���E���o��s�����w-_�H����/[���eK�Ă=������K�l��f�"����;�=�/��7��#��%��sÆ3T��կ|M�I�2Y�?�vl|��h��^�����.ן��;��C�3��Z�0MӬY*vA/�`�G�
��E��1l0\j�i�@#�D�ٹE��c�;�Tt��[��''��%��M�O�j}��~d59����r��=I�:��B�Z���9�0Eb*�k�u|�˱Vw;w�j=�);�}�;���;�mB�n1+Y��e>#i�L�i��y�^���hp�l��I���42����MV�������|Ϯ[+�ԅ$c�SckPl�ι��J�zTi�*�����~���gB�i4�z����R�J����F�է��c>���hn���.$<?BgW�@�o��*Xm�!h���~��{�����5�~ \x�e�=���ވx2a �p[H����~"�0O��M��o�U3:����燧�я}T}E����ɌQkg�G�����\}�52\��b����v����P�*+}!	'�iΗ*��\a�s^83��uwx��ŉ�u�Q��?�#EF���+�,<w�M�;�\->�y,&&2���{�V��a@f�M��J�oR��3��6�%#�|9��fH���~����w	�Ay�������.���OY]W�nS5��Im> o�?��k�����>�d�!}�5Vxd�sQ����Tj��]:��a!u����� X�&����6��=����Pُ��X�x%j.��w��j�Hb.�jE-�l������y ���S9r��`3�{�ԦB8{�g~�C��c� "ǯ\޶Ml��W�h�l��-t�x�3���sH��׼e�+�I�`����)[G�tkN�B�>��Q(�Jd�Ƈ�#aβ�k�0��b���jHz�:T&�`P��<�G�I�Ru/ ������NY�d������U�H��)?D�9���mu�n�P� ��/������C��q
΄2.��K"`�s(-M�Y��ņٺ�)�Yi�5����9�ߵÀ�	��VaBƜBz�z`c`�n�%%�O�h�t 
nj�DT��>���ჿ����;[�m�^��GG�������𢡄�7o��'��K�.�Ǯ��%v�$�tfa?A6������9.�����A��:+������/���F��v箷Î��e�W�¥��������cV	h�+�Xl6��֮=.l����c��%j��/�sx��a��V��?��}r�/�����=���|\x�]{�ĭ�0��;��O=N9�T�=�5��$�# ���!�)��|^�jEx��m����&{��J�uP|�-j���k�Z�Б=�����O<FȌu:G���V�wr�������;
Q��,��+���Q�|iH-,w�v>kstbH���ĠT�6)~,<��Z��CؗQ�1�~p?��NERo�ôK+Q�А����11�/�Y�~�m��^6;1���d�*�I}�w�5��d~`�����5��A��a�c�2�HW+ �.��g�NH���YpqѩɲG��ʜB`5��aAi-*�����6�ա�\e�uY�H�������ȷ6�6���b��7�B���/IMy�Ǵ��qBBb1)!L-�HW��(� �<� &6���GBA[�h���0�Uq/c��]�{��u�>���S��>������U��d�������ڄ:.�%�җ����*�/��bU��ť���c��?�q[�?�v��>�q=+��D���ʦ��#�3o������=�K"|xQH��DRL�yH�� �x�(k��_r�����wJ��q�
)���O>��"'Su���|F): p��	� ƽcRS6������PY����al}�gv�S��	Q���.9%�����d�	�����x?N�$U�q�y��W4��?�b�舞�w���#e��٤9	?k�9W�i �J���)hRE�bR�K����St�ۣ��.+ޝ�BT��zQX�x��4w �w��2N�!��L]?�<��{xw(��ˢ��8B��3��|�v؍鈕��8pk�w�g��3��U�C�l�sة��<�Ϛ�W�(}U���c�9V�T4�k�z�^����mf�X(s�x���o0'$K�M����{B�V6'�j�$w��ɵw�q��ew�˕L(6u�]���w���	o�M�~�6�n��a��X{�C4��K��Y�N�a>R��ׇ~��oct���S�]@!���B�Qk��Hp��P*��޽%w�3'��-*b1�!�T{/;v�lh�����%w�{�	�4�?�$��#m�ھ}[��ݡ�$|{�֋�Vd`ͫX'��b��~�-Q:�)�
MQ�����	d�(z ��=��u�ڵ�������9sf��p?t6����"BJpw��g�u���ND��s��f�#¸dѲ���KA�����/+��9�[{�*�q셌{+z�Zh��p5��p�\����{ �1��E�c֌=�N8��Lv�� |q�y෿��p�M�H���������^zV��=��S�|0�q�{���N���y��-Z�,lz�����k�f���nۼEψ-�5と5��}D�4%�^M�Z���V��w�C��ή0`kl�@�X�׌-��~�H���LSR1�x�����4��+��z�';�8����a�C�K��f���9��m�І� V��~V�ڣ�S̪����\�bad�Z��s�Mq�#*��0����6�TEx�8h�o2tj�ѫ�b����ی$�a��I)KE_%�w����F�m0�yO� �
w%�B$��T���vW'X2(xY�㪉3GZ���佪��D��.4��maV��C�p��yq}�7.��\���+�K�|���{��!�A����2���<�>Ͱu��'|d#��L���y����ԯPV�;y�B�I���u6`�a�Пz�i���.�۳a�<�c���q���?/ ��I�o`O�k��[�Hzi�`�e�-�n��8��@�y�Tqu�De�u��a��Q��^sM���,�����LL@q[�<�����ᶽ���/��g�I��t��^M��*�
XcL�H��.Hw��H�P��������G�yr�{߫*��n�� #�� �T���׵@ �zR�D]��ٟ���������ީ�c�c,1�|�{`|��@�P��"\���Y��8�U��d���{�x��}����GyDF�� T��|���"jʼn�-�ԗJDνO�C0L�J�Y�nx7,` ho��4;ِ8Ee�]�$�Z�T�򔾬�Ι�e ��
(NMM6R8k�=]�F#!1B����*[�!vq�s�*��.YD�[��f�|k��	���~Lg)R{8��#�l�NN�A�V�Y�*���_t�,���(J�q���b�l�4����]#��М��Y}aהw[A;-D��M����3)	����Fk���i\�)�ͼ���H<Ǫt(i3Y�!�L(�N���D�
-��m�(��DR��o����=�P2{<i����Wy������@B�h�� �{�%�HŧB&��T�4)���:9��S���	\��{�9�zD.�j6�J�0G�XT�*]؛y�h=�N��i�5ɹYS،Z>��-�c��Px�ð����^|A6��%E����yhU�ݖ-���K�xElS�%l߬��F8^�F&��7���s{�F !B�dѠ0��'���ر+l���"� @X�;���.�R��h>a`�������ۗ^��-1r�%��;n�-<���5 �3*�1v����M����@a����7�lT9�G#�)h>��6��XC�;H%@ �����)� 4-�����{�s�]g~C�_
P�Q�¹�:i�J�
������tR�e[c{v�T��;w��/�"|��o6y�R�����~{/�-�}t׎�A�^�l�itt<lyc��犣W��=��������7UL��Ƕ��g�ǳ�ا������K�Bʟ�˓5۾2d�uB�Z����/W�B��0����{l.�;9��괝p�ԉ+/�D��H'�*m9E;B�mA������t�l��U*%wE���Q��*�GK�&���)��J���[���FJͱ��3ޤ�2
iʨEN���sǝ+�ׄ�~'��xbD!�Q�����t.���˦�A�oٲ�5Ȁ65&i��s%=��ˇH9�Xo�żb���˹�;��%������Ť���ϋ��c"�e��0��-�l�^z��p�m�4�u�[�@@��[(�&��\��\��r���N�D� b�˨21�@e7 ���V��ͳI��G}T���G�E5�u*�<�1���f�HCfƻ���x~(���S��]�R^x�E��C�f�y�]t�x�H'!�M:hʀ��K������n%��(Qp1�Tݡ����2��+��R 7*���o��Z~�x���V[H��{��j��˯�<��7����`��
B�}�A� %�����Jn "��9�@���5�vV�ӝR༜��*�7W���]
xyl�a�Y���9 �R�����ۚc^tR�H3s-v}�*�J#�0&�L
�,rsV�qی�MN�3#�@�,NoYi.�M��s0�Ϛ�VS��LnZ��HGmFtι~�$�xXK�_v�b'�(���q���׺F=U��|��K�]�2�l mm����P/I��~T��!������_��<��1���=�>H�P�F)ؑ�5D��.9-�Y���̆ѪOJjF1Aw�oXU�w6�ټ(ڦ	��ClFKa�WvT-kѱ'��M�W�ɍ�4k��m�=�~ΓtkSt�}"IU*�ek�E{�'�"�yIPXCM���t� ؂��u�/�:ے�3��X4��4��:�Ͱ�s�l�!��Z��c�����ph���0gNoh�C����(8*��z!�o���h�|�8��r�ɲ��_ S�'��� X�&ō|���]�mm�B��[x���H1_x��H����(KvL���ʿ���	A��=�~���z�ٱ��(N+�a�e�����y�#�2�:�!����9X�d�p�	<����B�w¾�;`�9�/<��dOe�a���g>pN����'���/|A�06j���S���?���*�e>��vH������g������@l���N��g?���f�Q0�͜�jk)��X���f���;!c��'[��d���؂où\��]W2>��w��c��&����Shl�	Ɓ @3�]�\@Ait�vC���~n:�tᦺ��d79O��֌��8y�3��##c�����3i^�C@9�\ɋ/�[�J����CY�8ё�Q�U����"f�D�ٌ+ypU��&\��ެ�{K�7��0+@�J����)�jy�'DYƳ����r�BK�(d�0�j�z�[ SX����oCJ]�"�b�l8(����ˋ�V�JA��������<�T0��Y�-:��@�ZlD{@����$�s�G`�NE���]�;���6 ����(:f6����j	_��F���C��h�3H¦�����c�?���c!>��Sҧ��Wo �x�o^�=w�~���Yg���c�I���1 $��_~.|�s��f�zk�y�;�if�5�����
�v׽w�!����1o��oX�c����y{�z{e����H��f!���H1Η^z���E���NAU{�3�a��ژ�_�����������0T�rDDO6c�KՏ�PD�)H����%�D�`�1x����L#R	�HQ9����5��DP�z,��t�\�k?�ɖf�,�yG�:E4�C�pJ*������t����T�#��1��V�]m�80�0<^�*��(k�KU;������M*���F6r Sj��@@3X�!0��!sN�dft�������I���e�sUv�`ƫ���z}���I�V��6���sN�����2���7��3af�=E�?�9kQa�������D�����U��D1:��+�ƫ�j:��SQ��Ё|�]�\�`�*&�=_���ͱ�FFK�n.�U	o����"D�TS'�jԡt6E�.al� �T|�K���j���I��F:=�z@N�7'�h��Dрh$�Y��6,`�GP��9�U`��|�'�t�B�=2��9�����=��/l�ƺ�|���՘/�YKV�::\����~��;í�ޮ����GP|i�d��F�1���=xŊ��e���?�5��h��q�_��ƥ�\��q�S�=;Ⱦ7��5 n|��QH������טm<)jN�6d�
Y�+|ż�N�x���޿*�F�Al)�|x�W^y���d���y�Ў�vzp��8�o���������[��{�I'*���]L$�m,��믿� �@�Mdj���I}�,p	�@-������^�-�\�sO�͑Q�'�=�7s(v��k�
��J�o[+i&��ݢ���SMA�;@ކ6Q�ґ��]�eX8�����������ǔ0:��>�x����6At�h�+�ڏj�OUٜmGF�kM��Z���d��^ϊ(Ft:��E��	9��'52Ϗ\|���ʝ�&9Uѵ���Q��?�
�Qĺ��5�L�@�ꩇX	��J�3i�\%l�	�+�?N��tӰM<m����fRo��`@d�by=��sOTomm�!m�  �()id^8�B�&�0�=��
��k�;�$_Ң�_���W<�O]��L)0��/�J�1?���>)j����t� 
o~�5������H���<X�.���o�����N�
�$�ɋ���@��?�A}������Õ��X�/mzI����Z[E�
@]��<����� �|��N@�&%��=��߻Y`{�u1x��]v��&DC1�1-�6���c�嗷���OF�O��Ot.$p���a�m^)��ݑF!2��֓��c㍨\үJz�,Z6���w�Wu8z�'�,�q���JQ�!JDd��6�m]���(@���D��|��J�2gЀ�6�4w�l��Ӝ%�0&�zUs�� �]�5�{q^cN=��[�T8��_���1�ޤ���m�(������s��b����`<������j�h�w]�'ktH�����,�P��0@9S�1����I�:��k���/G���͈��"ʣ��lN� �����N�2�K:�$�"p�9�9��&�d��-�e�p�(�=7O�
�(����D���d�6�@��las�*��)�̲ާ�
I��o�a�4�Ai���杺��(z윞3���	D����f}�|����E�L��i1��G~FK?�\�\I�c��R1�@�5̺��b�z)��/�d�S�)~ �v��#�!�Xt�"��}���3LZx �;RP>О�Vj�;c\0�Z�]����>��U�x#��^X׹ȷǡ���L(=�@F�6�b"���ًs��1��s�j�
3t%l��zL��c_{��GE�JA��
[�MF�T2��{��T�M�1U�۶n�>��
@��z5�aӠ��~E��wJ:��#�w��k]�z~챇�ŅJ���3�+QPQ\�!����~W��k����W�#@MT�,�-�ܬ=�9�m�(q�˳���-�^ږs��Y�S�+m��[6oc��~B��T#�����o����(	�f�R�N=�,{�||01>�l���R4IΆ���2��d��/ޥ$�įoS!'�T�kjZ��*.���}s�KZu8T��
��(lV��+3e���e�TJ�`���5�V{�9�rn�wpm f�3n$v���`J��!�l$;�f�6)�@�Z��9zK5m�DK�&��}�aA����o�>��R��X��@���`�*���~��- �jd��T�,#��6nL^��L��	8U��0쭔2�Y��pU�oA�X��.].@�M<��BАf�R-��6-��xD���X�0�#BD���a�9��/�K�����&P��ٽ�--n*���M7����(a|�2O�g$��k�d���u�NR��W��^@����c	��R�i��  ���������u����������i�y�g���Vhɒ��V�=��on�p*2�?���
���N�=��w�U���6��Y�VP�|H$�Y%�HA�0<�?F�2�,��y������p�y��=��t��rک��Q�'�r���~�������\����,�i"�����/[.����(	,p�WR��ؿ�Ht���GQ�I4�Q�=��ߜ�K��ʜR��(�Nw#��ڼ��1�X��I��l&2^s��8- A�8�	$�y�������>H���ٲ�MUR�JW�E���dc�ao0�9��z���6g�Q��	P��b�U)u��������<�p0p�Rp��zP&�a1�zg<җ
kT��.���_8��F�Ǡb<���\r&�h�s�nN�
� ���N�����HG���2��sdT��4���=[����"Sl<�;�0�{P$�8+=�'魮�b߷9Ƽ��8{9�B�R��74=��&8b'�����L.ʌ�D�W1j)��~��R)�벒T���ǎI�Y��
YF�/���UxG��|�;�b�ͻ�˞$�b�`�y��6�(�{�Y9X�$
?�êUkd�A E8ù�QF�f��Tpǅ{c�!k�  �h��{��		hA�Ѥ^�s�㝊XP��փ�E�{O��Y�RE.�Ҁ%�8�`8� ?���dx��gC��"lz���9�`�v���Rf��cD<��2�����Wu���v#���B/�a��I�����6o~8餓��m���sKD�g�ȕ,�ҥ��+���tP�&��wݥ�MP�����s������
�\ri�����@�A���;5�W�_�����46���h��oVb�>,g�TD�K�2�I�����^s���������]7wlxL�����k��1ʆF=ץ�/�N��� $��C����~ܲ�b��K�r�R �R���au�3N���P�3�ͬ�S]����n6ۼ]�a0::���7*�d]�� yB��������[A�����);T!�� �}cS�����k�d�G��"��Eˀ8` ����$���M �DX��t2��3}S�Ya�Gx�
K^��g�:/E4*Go)�%��H�AuN�������dĝ㥂�Y��4�9�عC/o�!s�TB�L�Y=]z!���p�7n�����{������!��ԥ[TP���?����3�ٰ� ���o��o�C�.�C��!�Ft�h�R3\�I�ۨD�Ic�e�Hj�`<i���b�-ѤT-}�Ea���^��s���/�R�R����)Ê0cFZ����9��ׯ�{��b�.}�I+����+@��K�/c:��F3z@!`n	��+���rG���L�P�w�ĨL���80<$���=�������=�_ wDz�"��R��$��U�.)��%�B��F��fN�g��tQٖ�6ʖ�c-���Y�'+u!��p濥X����c5*�{�F�u�"��y��!�������ã«�(�9������U!����Ÿw6��M[,!��F��ZRa˯s�"��Ӟ�jl\],�ķ���z �E 2���ݎ�a�t���>����Ae6�'�~�L6vr�ȡ�������G<�����Hf�qD�-:��i�lS��j �S�<��U� }H"su"��~˪9��>�9��*�٪-GY���Y"ձTeS\��r%&zF�߂�;�0"pT@� �Ú�pZO6�6b.�Q��þ)�dϑ�����G��'�ɝ0e��k�k��8�;���Q���꩟k� <�a��.�<��~�4@2:�]W ���Ņ34ŗ9Ȁ�b?;��;�
2�?�8�D� ��fY�O?�L��{�yO#��=��?�H�}��ڗ��7�t��,����<[�'�%��4�"l,��r:�_�1���Y�q�h���~��)@���$��L�4�ن�ſ��y�g���Q����Ƚ�
޻�裗˶�M�Z�?Sz���=��hC�%��x�ȹQ��^佨g��v����P��W� �Fx�8"��]��Aյ�ڶLb��'b�@a;^�ya�TOf�#�_�$Ͷ9��Rᤊ�"����9ة�'�^CD���3{��Vw�C'�^���|��N�@�����~�t8��SO�l,ޛ�X��S��Z�R��d��ɠ[��P��.�ރ��"��|Y/H�qȝSͨ_��Tv"�C9#��L�G������E�W�
$���lO,�/�ɘ�a�~����F��L��KoUr��Zl�l��s<�d^�0^FO�,E��ӷm��(�4@y����r�)V��b�h�ؽ{@�����l`�b�+���Ν;;����x��[��:D v�vv+�L�k��&cݰMP&��:��,�Ȯ^�J<�Ո.�]�#�g����/���ѱ�X�xcL��ڵ �p;N��T�QY�yz�}�b��Dv��A�Z �Q�8\���ɶ`��� ���i���(�۵�eT0V���4d�^|q�G_m�~��h�'��Õ�|�$g���4��x��0/0м{�1�6Lx�P��+�د;���n�g� =���*s�M���P���|C~�E�,
sN��J�ю�λ#M$�¹�؄���#�z���ݣ�M��9'�� �1_�I �p���T��b5V���^�=�V�*������g����Ɨ�o��8��Y�D	�Ek1��c"��(;��+�E���gp�2�#h-��A�*\=Ġ�3��]A\��?���ޫڣz���_0Wg �쌯g~E�ȳӑ:t����ʄ�w�5�[ۣXR{���N�ݤ؍�b~2�[Z<]�rH��U� ��#��\�11 �'ŜQ����|��	�Mvݲ�}l{p�[�e��M#�N��ʲ�1�jC.����0lv:9>	�9u�b��x�ѻVc�1�k;BA	��ew�U��kU]/�>�ZgH]�<}�+*Qxt����+�g��@uP�	�99� ɖ6�2ѳ^�6
�3bA�cV��jMh �&k�1�3���Q�����ma�ఀ�ˉ'�N:q�w���]�����;�QG�z���6���ʼ�_Q��g ��YH!�98����4@�/�(Gw�֭�J���ػ�;\vp`�$7�/_���.���r@�m��\p���ޅ�$P����{t�T����{ro�?�J ��kd�(r��R�@oB:�Q�ϗ_~�dw�(�}>�g΋���Gk�9�S����|?��p�"���{ w���Ը�	 o=
Z���*� �![666 ��v�gm[�mU��9�-�;U�84_���}��c��e,}�JIT 9�Eb�w>�p��k)�ηM� ����@E�ЩhP��$����q�S��h8!�B�1��&d2G�y�aM��ˊ����9���u�?��kZ�� ���J�F�Ź�SIUZ@�Y��,]�X�+��\䷤^ռ����/g�M���=��&^��p�����)����&���w	������<��gfu�J*L;�P�����6-�yZЕr�#���)���#?�d[�D�9��b׎�p�Wɣ�ַ�����y- �=�F���SJ�����\�� i�����?��RLf�|DC�ay�/zo��CK"���{�N�(��ٸi����C6H�����a0<�)�ݣ�Kg�u�z��|Dߡ��l-`�w>����ʳ$j�aaC`���%�NOq���[@4Ɨ{fl�J�~�ế����7�Utn�K:�@���H���⡪p��ޘ �����=�:�护�Q��E,cn�`���)D	��XI�&�ѹ�p��Q�JE9��c���(�]hu�O�׉�
QT9��l�c�O�f��~���F�&��X!z���������A/�p������6�Ϩ>�������9���HJ�n7�rÀ���\��o����Z�!�
����z\
�f�����R��Q8�;&�e�Q���1�! mS�I��"6�E*�+!WVSp۰�nR!�\�>z�W�8}�m~��s^�'�K� ��f��AӀ�|	`�o�a�]*ͣ��p�ژ�{LNNE��K�T��]�*�R�׊RU�g��V�S��d-�/����ض��s)�`��Ȱ��(ѣm�67�H���c60٤����8֜�K����l��'����H��;��0k�<�t����p��>�̳�����-:o�3�dR�MfgS)����}4lzi�Ҕd\���3�%4f��b�Pe��ZLGΛ�E��?R�B��T_8ͬ%hAD��=��ڳؗ�h�ᄂ�+ڗ9�8�\���Y �P�~��裏iL%g�!-�̮3j������a��;�\p���A'�����la��b���e�<�U�{�E�_%�̸�)�ٶmD���t�6��Os� ``O��I�-��B@۲e�4�{�9��#� )4䝰�1n�c)�G�D�R���(/(Y�t�>ŉlW��,]�OKp����Dy�c����(dl=U�?�3�����ã���Q���Ƶ������������l��Ml�q�\Fb� /��n��BYl0���E�f�Jp�R�hQM�e�	�P���l-V��&uCsl�Cu�ѥB�o�B��D^Ơ$)�V7j*�$�"�����o�%.��@l�׷�
�MW��z�D$�R��l���ڲ5��;(br[����V�hf�յT���q���ǬQ;#�qN�m�ѐNLy����[o{{�k����~��w�uO��_'��:QF��p
��P�*���J����~)�ﱅ����o};�s�٪:k�kg����kJKc<�a�q���}��e���^�觪�l��1H�J��:1����?�f�>���xU��wɀ���
��x��U*�a��2S�`���������3Os��=)�!-����1���/����l,/�𼪺��8������n����K_�R8��sԍa����n߸��q 4d�ms��J�yj6')nb�@J���/?Z��0��B/�R��E柷�����y��)�(n���b��QT%H�\N�'��Q�ʿ�fH Vs����{���F�*�)�[Ez�J��yT��=���͸S%�y�� &u��6'�]��$�2��8p�'�ġ��/�pD��T��W��dx!0��T�ȧ��͊��RtV��2����t�W�e"�,S�(TK�j>��*W�,���R�,I��玢�!̨�V�^b�8�3
Sشs��(s��dj/X?,��>�C���d�ꑼ���v���A	jW
�،���Iʳ�(��>�=K
-�W�<�&s�LKC#�1��94���9��Q���Bg��P�1���j��IܒT�K�Hբ^Rזf�pH�h�G�i�O�W+ �r�ߴgPһu)���<� �D� $��1�Tm�x�B�!�J�;ڔz'�**���lб�&ğ���z�����-atlX�����Rᣁ���6�T��C]�}ۙ��Wp��g�3�(~���}�����N^�z^�*�i�|��޶C���B����a��;���Ć��G%y�3����pض���7wA8��^c+��A���?�Q���YڃT�a��'�V
xՊբʌ�O���L��O�Acó�}jM�>�c������h{ª���6����Z>��?���6�Ͻа�2.[�"L��VIT�
�`B�����d��gJ�^� 6�����&@ K1'c�� �DQ������]^|�Y�?J�C&;�t�Z[�����k�������|���i`�4�.��{9��j�K��V$߈��-����YբH|�*!�F��}��y�F�k����'�5���*&�k�ź�Fe{��h[�D�X�Z��Ёa�+�<9R^�9��P#����֘㻆��(}9oh�h���=������M�F,�ȡ�wH�j�"���Gų
!9�6���}i!4�2�\׋h6�[2�H�#P*Mxk �h��ͪ.����>SZ,����)�4=�*��xW�5\�T��ш��C�KJ�qM�� ���C��v��+f��p0X�4I)��W��0���,*f1pࣔC�]9��'����u�[VQ�իׄ;n�#�r��J�Y�>�9���=����5���L���?�<��S�%� �����٨���u�N�gB�U�-��	�i;ώ� ���r�3@ }ʞ�7}S�:��Եf0�Hb|�!��{gA{W�6��t(���q� ��NU�|�@�w�dB�Y��1���<P��uh���W��s��w�X�
��Q+W�@�Jo�Kq�ڵkC����6v�����
l��&��{�Hs�gSk�];dI�/i_*�q��I+'�l�WQh�F���w���&ݶٳ�F�v������[���KMM�|��H���#�f���Q�.��9?ͅ���@���v6z���w��7��ߋ��Z��6%v}H26���%���8Ҙeb�@Y�(�R�z!]V�e^����o�j1P�Z~����,S5_��?t�G�oL��DO����O�[�H5��Z�y���c�wnS(暴9��&��k��]�9IJ�f�QE���"�f��4��V-�;l^�܊9��L�ژ��/Q�`�a�љ�d/��I|]:�f�I�%�R*f���
qߙ�G���(cQ�`�98c�(�Ӣh#�B��d^�A���SH�������j��c�M��)&ϑ�#�М�TL)�!<��K��-��ʥZ��)H�1"`���L�H��K�@:�H�܀�����iD_|i���A�D��Hq�dI �s�/�"�Q��dW�.\"�[o�U{��FH�}�s��9�<���=����̓뺮s�}' 3p��HI�H��l��d;��<�Y�s�T�~��t�T�^^�{�\�_&;��$nO�H��Y�cM�HͲj$)�3H Č�;��}k�K���8��>*p������Z�[�:y�ە���^�Ēz(-]�X6��%��=H�'_h��#ɿy�w��}��_�u_a �����ƻ�;j���S�(Ɗ���5���Pa���sy6\ş
�Ȕ����X�2�\�,<���0�`����۟��,T���E��D\���en����y J)[�W{V�1�g�/zG��S'=�Q��N���F������-w����S-�-������Hk��Q$>������p����.EqT�L�8|(��X���>�z�H_nM��7�(mL"E�(j�U�K�D!W�-ggT��l��Ao���юDJg0 �2@�D�Q�%sʱ�;yF~é=P�{�iq&-a��!d2�̴٤L���X�ͳ⺇D�XD���퓠4�� &b�f�z��#�P7Ư<� &x+6o=w��qq��]t��������y�t�\�X��n@	>: Ѧ�63����� ,=j�d�O~�Sf엄I�ة�c��_$���ވ�)�7�F'驽�#�1��^(F��YH�&�/^ ��Y#
����b�b�1����?�l ������9�+�;D�rm�729���+�)���ϑ��9��<?|�����N<N�^����������M�Jϐ�����&^+�R �x���:z]�v� %M���S�( 6�N,]�\Uy�م2p��1���2s	#�x}N��(=��x�]]����W��5Ϩ����u�%��<R�/�Ԣn]^OR3��&8OR.���� �Q3�.ަQ-����5>���*�Epl�5'n���*�Y�4���Job��F�6$u�w�[���J�ܹٙ s.t��j%���\ �1n�J��j7^�Z؀b�NZ���-��ؚ��8����M
��l]��'Bq_�Sł�aa���M�f��=9�z�;7s&��3�L)�x���3��DF���A� �151W�/8�0m��G��A
��YZ�Ě/I�/U��Gm�l�E��)>����K¦K/U6
i-�QT�.Y8 ۇ��)l�Q�J���<۠M�۽K�גH����UW�V[{ػ�^{U�`I9�ڝw�>���r/[*u�1�ID���]j{�Z�v��o�x�%W-��X�Pt�C��\�ג���{��������Wd���+;v�`�R�Q����%!
���|��`#I�s��W02~�IA���罊�? �� ����+1l�{=��S
PIg�����H&+V @��#�*Gd���[��V�KJ�����?Wc�L����<��
暿��o��{4,��QJ�������W_��+J5�Z��޳@Qd*�-U�z�?�thkm��[n�]A��_|I���(=���v֜mh@�8��n_�@��d��J�u9R�z��3�! ���G=I�и��<�L�ޞ����g\j�#aH����_�=:bc�o��94]h>��&+����~���u�q���v�J+�IC��٩��y���a��	�U�q�D�ք�]�x��>��A��5�]3Q^~�SI6 �QG�X`A#=�$%�G4��0�����i���3h�p˦9;[k̐�%�w���v�P2���h���p0��h� �ȑ����Q�2�^�f��A2��mrK�2vHa�?h�����X�Q�5�X�I)��I/ʮ���M��H���� _�fMȣOV��2��10��N���K4��o~��� T�+X����9�il�, �J�� u��ŋ� 0����Ϫ�sah���X�ͳ"��g~������9�a׮�����Š dyD%1��N�w�'p|�����}�cw��f�6��Y�=��ZԇuB4��S�tƇk�������N��g�f��"�� ��� ��
�3���p�r��@k�k'��a�E��4镓I�4�l��0Ù�G"�D�kQ�!����ũ�4����m�զ�d<HG���ŵ��F5��>�mE?g3��2_������F�?��")��z���
ˈ�Y�Ւ��Y����J�F�c6�L��Y�W�s����%�֕�G���1�~n�웳'�~������u�8.UE��ыY�%�l-��҆>!ii��&a���t�D�i�-��ׁ���ix}ٚ��(��z�P�Q��	2�v.m�z.�2f{;�Mb�6��ё�ӻJk����r`D] |9��%uZi��J��"��na��Ȱ���X#8?�[$�@�p��E����~lϜ"9^G1�p��5�pel� )��z�I��<<,]]�r Y���l`_�g�d|*�ށ�>�W�XjcWD�p��l�d�� 6��@��"z�k����wܡ��h�d���>>��s�!��{c��}6�dN�c����s�]���� g�<�����xb�ٯ:�]�߻S�dg%:o�����`а?KZ�^K��n�3q�߶M�*"��Kx� X�VQLJ`���=�y���p����g�߳Gc�y�&e���կ��9~�M�s� ���g?���>p�{����k`h��u���{���v�XL�5+K7���u��r���g�3���/�K7^m�$Z�d �R6��.�dϪs]����%*F�yK���v���zo>x�����3�E	K��;q��L�[K��sD�?����
h�o-kk��Řm}����j2�����QD����x�ة�>6Q�J�5�9��Q�j�*��6����-���Tp�	Ah�n��/8љ�J.l�����i��A`1��7����=]����Iq&�M§��	�>��` �-qc���@5�x�<B�_��W���x[5���b�s.6}2�47^���t��Ky)<��s"7stv��\G�T�^�#Ǽ��<  ��Do৞zR"���o��-����P�IWL�UC7C3
mv?D�$ň�N����Pœ$5{�EI���~����3��C� I�@��t��S��E�h���d�&T����+��]���Z�pP$(GB3s�Pp  ��k��wIE����?�0 E�	��VS{�>"b/��Dpo�7�0�⥋���o�N;9y�T�qn6#o���%��&
�T/r�����7�}Xi��^U==&�<j-�a)6"��j$�s/�މ��1��vd�����߳��Bã�K���j�z�P���Ibe�p�:T�#4$~L!�9_Q�����ZQ�"x�$6҂-m6��T��<d�a���Щ��)�#F��D�Z�!���>�&]���n��M_�����tp���=WT�&�SU��r�΁0INdԖ+ޭ��	)?'Y��Қ�r������i�l����pQ�9�H�ekbEts���$�t4���ڐ{I�37v��{���w�#��iƾfk(�9g޶����Zۡ�ؽ؜곿���AƬ���ʨ�PE�G]fO	3�kt=��ޞ���۩T�Ωm�=�L�M��'�W��cUb�-��ƈ`����*C'sS�ؼ�*9�7��'ϼMJl��{FN�gE�C�=���OK��*;wy���BV�hܼY)e�Xd��-NN�`箝���8�)H`*N �m� p��q�)'¢eK�SD��H�m��q!k1��7n�V*�*����׆�����H�	�L���5c��n�V}�w�x�/����emC!J�� ?�6[-	[����?�kA�[�سwO8b�&��S'��K�xY�ȅ���l�T�O֮^#9��� X"P�$�ɀ:�`������Fi��\'��)�Y����*�v���a��@���k��X7d���H ����p˟y��pĞ����wQp�=Vj|�9&\:���Gl��^]�l��e8�և�����8�-D��� �'%%����̔W#�gv1#Lѥ������X0u� �.Q������)|�Ɂ}�dc��B�Ⱥ6jv=�o�a��n��h�c�N�2�Y�zEEj ]�lj[̑��U��sr�����Ტ�U��1�nj=��TA&��l�J#��Q�W^�M�v@�8��m��$T�2n6�6%�X�����6�,��.*��$`=�P��z��1 �t�U���Iz��	�>��&'-ya���F�Sj��z���c�	^��O���� y�f�W����H�֭[�3�"t���ݼ>�M�KZ��_����Z�>��'��'m��bB�峟��&�����E#��`������l�#���0<�����i���r���җ�$*����OJ�L���&�3|�J�v�0�:O���,�A�	/�����Q�B ���	X� l���3���Z�.�L�����˿�KI7` 0^;^y���J��H.�l�y��u��5 �`�9�E�K�hR��?��h��e���\0�DQI��X�B|����&8�ʶwx�ϡ��Gs�� ���{� <b �j��F��{*!V3'�}��8mVZG�6NjN&��χ	���3)E�T�g�m&F�I[dő9=�x��N$�g��4	�������v�1���V}'N�f6k����erٳ<�������>���#]��1����w���q6f,ґx˩�'��Y�J�*J�ȇܝ-gC�%����Jic%���\s��|%�t�g��������w��t4�ڦ0(o�W ݕ��03:���LtƉ@R��3�W���NP0�<�x �F���yH��u�4 ��Z��dpm ��)��F��ᑣ�f���6��KQ8�0-�9���w-M�ĳJ�Q���b��Ǡ��Flz#���k�X��\��HFlK҂�TJ1�W՚`��޺�\E:�=��	�@��EE0�/���0�O�毭m�Y+ g���R֩L��y�%K��T����Ͽ���ᇢ�=�}���X��g��g4֮]���Z9��[(>�5�-�>�m4�!�,K%��;)�0�^�~���.)��3�`;��)��Z򼰗8� �n�^���Bj�1a��E��S��s�}�ֲp:(;�ћ�."{4��^{E�kp��;>��k��*DlG�s!uM�k���g�|y��-T~{W��h^�t�S��m~�yK_�S(��Z���xL���#<I�w��ϟ㕍T6
-���:F�;MOO(��}"����(
�sj�73SV`&uK����z:][�>σ}�%yr���]-^ˮ�i2�o-�s5$�_�:ھ��ו������ֻ0}a��-~�(5&<����r��-�>ݜ]8����ab|Z����^�H�D��#�|��ضo:���G�V,(�7|ԥ8\�7+�x��KB�iS�gR�It�7U�I�-5�&dOʁ��C��J�6��X��U��l��@��-F_8(�����c��h�j�=�b�?!�y�\��9w	��֝�Bi�d���S͊ի�.��(H%�����׷U�!����N/��������=qF������n�YB��W�o����Q���d}�ӟ	�X�E�����J��>�
O�ҹ	�p���牑��|���3v�zS�%�^}u��mI{�2���>�{������((��z��������W��F_�P�cl E��Q���w"�_Z~�CV�*�8hȵ�똗��Bu����uQU{�����B�o��~�uq���r��+������K*� �J컛�@jWɦ��2�.�1� �㺆yq"�������|�2������ ��꬀x=�i,���{�݇r���b�}��}H�(G�(<�l�\p�j���8��� '~�%��Xލ,M� � �wv���U*�����z�4��ԛX�� ���z�:�J�_.��Ѹ�w��/=�NY�]��3S�����?dg&Ci�t(M���8U�|�����Z�m^���#*b�^8��1�/y��F[�U!�f����KV��B�L]KY��\�\HǢ�hA��	�Ej�T����lCp>5t�ЦԤ��!٩��4y��LA��?�o���C
p�,D��������E��U�b{����Da�O���L7�86�p�wؼ�쳖���z
���I�{�s^}y)2��C
S##��˯�����>��ңݽ=a�}:,2�*���������v��tR5�o�z�@v��������¶�k�0�}����x[�v�(<T]c��?W���B����ڠ���QF�U����H��HF��q4{ �D��㹰�$ �I����I�c�SIt��4qK9�Z�l>��{����j`�-I�1x��/#�Gî��¢���kc�u$������.X�:\|��06|�lnVω���є�)�=u�P��"���ptxFD=���6��|o	ܥL�l,���b��P��c�����L�&P߆��q�7cǳe��_H� �%	Bdk�����(�S���Hi�dhd� �c�0�f९�s��6��21*�f�U:��]D��ȍ�6��� ����k CH���ѦDUb�P�����M��jmޗ6U}�hD�BLC�E�?�J�+o�5��㷬�ě.�4l30�ԞF[�`�@(�/�ځ�8��,7�6i��>���AV�uy��)������ժ(�W1ˢe���Щ��ۧ�mp�6m��k��'��M[��[n�U��x����S4�t/iU��x� Y�Q��Є��ޏ��N�R�$����)��n�M���C�K-������H1�E9΅���2�I�2� x(�)p��� �"�dƂ�"\���������&���3�3��잉~�caU{��)f!*���x�U]��;��W^y�@"��2�����ydc|xxT��N��C�ޥpkHc@�9������ѵn����r���M�`�b8����d����+s�_^G�ϒ�����AZ�q>9v�!N���xġ�T�%c�?��3�ל�����Ƌ�b����l���)�R��w�U� ��s�x7��?E��X�-5x�鼤�I�f�Q˕N,�J�b���3����b�!7�A�lG�E��wޓ������v�d�d�Rt5+=ºZ�a�f����C[�@���4��"<�\]�&r@SDCk�P{8N�VA
Z�5fH�ĉ2�����N�o"	�b�5c�	ՠ�R�Ѫ�
u��E���M�x���+����F�W�d]Gp~�=Z��f�g�ٲ+.�\f�4�4�6W�1�p�YX��Oim�23��E4i�lĊ�ê�+\�jbR�f�bAN֤hN.�U���R���fZ��Qzܩ$˕�*�M4���?�e~�;ߕ�6�f��o�̹���Q$��ϧ���'�>$k���F�`)rſ��d�(�ys����ޏ� ����X���6۝�Sp�aT�A!6�)�v����gN�d��M� �Zx�-��3��[�u��m�l�{��o̠G6Ŋ��q�/�=���/�2[��}"�Ƶh��w��VN{�����G�HnmE*�I�ck��r��t?۶ݮk2L�ct`����~��?,^�H�=hC�VQञGgwW��������+�')�T*��eOf��3ب�q;'�P@"?����L��-�h|
�5ےT ,���	�𣦂�%Y��
ᄦSw��4B�D�c?������|����n�0�@�G\�((�Uv!Y����'G�Ck���\K�АwikoW*��M"�dW�Y�N ��h�����W]uE���)�4�-�DZ�l��E�O��
$fRg�c�~pC�(f U7`�	|�~�.:&���8����z�R}KԬ��Q}��p��[�Q�;l����/;�Zº�1Zh^ƴ���G�'�7^p�>�BJ_�%yݭvmG��]��[������?|ߍ7�{8h��Ƕ��|*}���Qy*�2��6n,L"� *���7_��ۿ��LÄ"Ō�ǵ|�C`�ϡ�L|�a�� �{�}��[���Џ�`x��W�w�)����j/E�6�$���9 �[o��Ap�B��p@ 1oD��H�����~H�|Fў���m�&�0�&3����o�r�"���}{]�V�y�$7�ꫯk��i� ��k��mٺE�Fn��=a�޺�UG[������ִ�(��U��j���n�yi��=aH���v�|� ���Sr Z˘3�AT���Ȑ�#�e��`���y�"�g��������`�M�%@�,�R$��"��=h(��z?�N�Md�I����^uZW��>����"�ƞ♳�s��2�(���Vѿ���4u����r6M�KA��{���FKH�Y�Ν��R�sȃl�14 '.�Ti�e��l|~*������b\Ƙ�o��WO����#�g��S���k*kS_�\���N�l�;c/����E8��G}�J��l1T
3�m�Sc���3�U��q�
�Z;=RH��� ə����U΅���Eng�Z��=6o�v�<.Z�X��\�#F�rڈS�H�\��@������ry�5|��|������Wk�b�!gBZ�bƖ����+��LN�Ӷf�����钂Ls�(�F��8�D)�G��*]+���`��gyF��֖�������p���ߕ���h�!>4t�eK�k����϶=.
��٬G�����\�r���Jt�0�|̮u̮;cF��{�2_��N��PÁ�f�(c�.7�E��If���M�٩B,���.r0����a�ɸyk�	��3�5�Q���=D`�����^q��RA���'*��ę���(��>��H�8����.<����ѻ�m%bP��'?%�)v{F��s�ݻG�~�k��*=L��FIg�8�P��rK��+�Y�cP��Rw��-��buB9��@8|p��s]�&<|����e<��(��mQ��� �Kv� <P] �?�2��oU��	���(��|Xb�G�
��������+%�$eSs����*2-*Z�ݰ�:C�Qg���|&X	<���;�>8�S��p��U���|^��8 N��&����PɌ!�4���Vzq^%��ÿsQ�-�`c�� +�D���}��Im���H����x
��9<~Mx�g]�"F$����k�.]��l�B�	�s���xXxQvM�D[�|5H�H�����Uf�z ��x�d5x�,�j�k�P�oOק2����u*|�?P�|�.&�O�w��7�����������`���\*����A���0�K��}$R�\�E������t��r�?m�$=d㊜ ����g#f�[�i�*�̸^r�%�" ~��-J f�/���p�m�kƠ�uI�@d�wf����p��/h���R���3O+* � ���& ���أ�)��&��N��ďTo�B�+�hE����O8Ix�}�}Z�pS;�C�� �ϑ�%]4�B���.��|�x;0�t��?�j�ב�`���f�����A[�]t�~�V�����l�6�����T/�����f
�4�Ͱ�>yB� o��O�b�E�.z%��D�#��p�_�� s�B�E�^潼��C��q:�ֆ��b�9��U�B4�Y�'��8�w�Q�sV��L�� ��}f����%��c��|�8<z�=���/?R�p�W]O5v㉟g����#������Y-�u����l��#��c�b�(m�z�G���F�{v�:���)+�=^c����1[�+-	��k)"��^S��5Z�bK��_��W�{S�����X��6�ӓ�(������q��5�������
S��a��ʸ N�S:�ִRȶ1� sty���1 ��%RF�K� �H-�Ec��j��0`���_ ��?�B<(=����quiaÆc~���Y/X}�f�,�w��-�e���I,��J�:{]E�,Y�(a�v���Sȁî��������~F�i>���/XAM�=Kc�Q8��YS0�ˣ^D=y~˖.U��0��K/��-��}H���"����k�Ⱥ=��#jO�������'�?��������L�:��\sG��ꩧ�ўy������Zs�;��vi<Z��e�g��)熠x�\��={��2��[�z��b8��x�w+S�  ��IDAT��G��736�Y;s�Q2��������Rjڮ��:�_��D]c}Vcf�Rq��\����C���,�gH�}F����̵h�v%�&����޸�%.{�� �x���̠9q`��h��jsh���d[�sȸ��0�h|��B�Ů0�d�d0�����E>26*�-=�0'á���z0�Ql�<��vg���7C�������U��'�FSQ
�-	h#�I�
��1��T�љT����1<���N#�������\�O���w�a��!V�[+0(��da�$�c����{�<%$��+|O ����C� ֮_>���{I�9D�Л"�`�Y��O}J����¶��5 ,�dr��u�k{"<`��(������&UW��U�����0t�G�
m�lD^h�}C��`��f0`Pe\<%Q�57<�e�.[bcqLw����߾W���^}C��1GD���^jRi�'�خڀ+���CU^�c84\+���ȡ!ZJ��JgfRj�]�4��(����P�r��׮]+���ᒴ�.�`�W-G邎�b�������T�e����=zH�g*̆N+E1#��S�믷���o�6�/�j�$ĭ�(�����.��&����]��ɵ,Y�H=�-�O2�3gb,�f�R����ɣ��Y3��ҵH�*�����k�g����h��=��Ql���9��X,����ezrg��CU���G��D��mՂD�X��l��_Ql\i������%Ǚ�LHg�7��XLR�D���\DX"��9@�:�d���:��-�������W��"Pd�Wā��3���g��S�c�w"���5K�adjB�3��G�0O*,��M���8+転���žA���j�(zoO��p(��S�>���'�O�4Ȟt�������f��S�����=dN����8�����T�ZG� [����P������V)�}I�o��Z�]�(���5�<.0��l՚p�e���lݢ~�tH�[6B]�b�	 �Bt�ϸ�+�bG�����6�Q�y�U�՜���[�̳�([������6�H�t<��ԅ
���j�'i/ġOZ��7_�����BE�i�	b�O�X�Lmm��`�Ʋg������-��\��, s &ǃ�(�p��AM�:<G�=�?�'���������"k�͐E"���n�~��=p�[{�9	�h_�ne��/_�H{��Ͻ�^��Uh-
l���N{W�b�w���$�ϔR'�EAQ-j覴q
*�ǔ�g}&��89���z��B9
�;-�k7���rI���HgU���A%	��Z�ϙ�������ͥ�\x_��\�3�-�����Cm�`l�2�V��a���"4\�z{%A��=W@�d�(���i����#��Q��l����Ԛ�&!c	Jg2"~�Phk��;9<��h[��7=�D�o�;�՜���W�G�����Kz��D�	��<@�,"�.=�R�8�ݘ�T���$0��N�+��ZE^��i	�C&ϧ�G@Ba����{>����֖i�VWl�n�}���L��T]{�u��F|q��s��yX|"� <��Y��Ǘ�,����:���Ǭ��=K��5��o�W��X,�(視���)D���Lz�C!yĉcSq!�����%� �"^}Ay.�l�A���&t��O~�E��7Qd� ג��Y��W�������]�qЌ�ظ/T6Y�Ud�IHJ���pT5IOf*����8ׄ�9����H�M
Ǐ�����kք6�s�d@�,�e��Ih�!-Q{=�����xxZ�*�W����r����l��!Y��C�e�P�k�C��+� ��8U��I6�.�c�8`8⽔�>�̻n��v&����h2g��!1��9pt����{6� a�cO�Юy�PNM!B�@3���<~^�����֘�f��Lx�C�D��$)TkA�d^c�7�JVQH�es��-���s�ޟk�q�8M r�Q��,SN���6gm�n�u
�,՜bPV��9	&�rRHri���<�>�޲�tuk�~�*Ԣ��9���D�"�%@��Ϯ.�κ"m�#�K<B�Z�9f>`��V��蟸�|_����-K"��k�C=�����e�~�1{kϛf7���\�6�7��#�l�b��7p0�����۵{�7��qx���ŏO������q� d���`u0����TȆ��}�2`I����4�*N��X�Y���)�G�6_� vm�x���P��=EU���������>vpEs��]�q���^�(_`���0���ŧV��\�S�J�^�;�|����*z���{'�w��`x�7+�H�lҒ��R���LM���#�.�s�>����j{.`�#���*�������Q���J����j�H��T�<�&SUty��}ݟ)�	H�M<Ke�bFV4#�fj���J���IsY�߼�H�);'ǥh���t�S����P�V�����m��v����� #���X�7{��~LM����D���ل��I�n��݊V�lQd�ހ�\s��4(�����cD7m�V�ЄCz(��X��U=
Wi��������7�'
�P� �X8)�����%D�\���#(]��Yh����Tl;�sV�.m!?�R
,x
X �a�MJ/��B����2"x2<&��I��޽.����3��{���=���v;������a�@�`BJ��������D�x����w��Ġ0o��j�����>��{u��'�c{��?�|����7�d )&��1��N'xf�NcםZn������%��7��L����Ҝk/:P'���)��7�N�A"BH52��j�&�]�]~�{�s�ӱ�7�I�$�Q�-�
�Eh#�M�f��mZ����'E r�c�3��Pmm�}��XpT'�A��'���jҮk���Â;t��*�I�X�2\����K��"���o��C4D��k�aT9���ƨ3������6��6����0�9��u�F�_��u,GQ\+��ll�I�U�us<ZU\'}g���N����9HP�ϵv58t�a��ΓRN)��^��3�a��4��<�9�Q�7��~ެnsZY2^�ke/��sUffì�|C�s�����dj^M�V{�@s��k�b����X��P�9_a����[���1�]wrb����m����E��N�W�'��$��9��k&#��wD�՜���Ѱ~	�նyd(viQ�?�Ü�ϾY�I�Vw�Dn38m������q���F���lhk�T%~�vG�t$�
�8>堥�өzf�C2Z���H�V��j������ ��j_���s@���";�DY6N
���Z;W��9z��$N'�Fo��N)�X '�ZsY�ɱ�pBZ����աԺ�>g'��<,����'���w�����!Y�qg�:zz<<���a��5ᓟ��l�&
S[U�'��[�%���O	��ʫҐ%��07��g�����@ ��DϠ�t�w(s�w�^  ��B�L�\�m�2�~�6�HĦ���=y챟ˆ~�,f<y&������d^���V��?44hέg�o�Ϲ'��UWmQKU�4�x�e����o��7y�!N���^e6�4�����5no����,�yc:k�gc�%k>��	f����}�U�Q�2-	]6�$3e��FS4}��ښ�)��? L��͹?iCS�[s�y�ñ�u)�+�^X�7��^]'�B�Y���4E��뻚z@�2p+ǻ�Q ��9�-'�Ka�Ƃ���A�-�%vM��b�(&�_�����-V���Q�B����6�OC5d��(_���_����� �B�����T�]h�62��˥Ơz��ՈDOH�u�FW�2\<;3���7_�Yag�#"r���V{)j	� �{�u�k;�`W�.�D�`��õI�'rRoi@"��e��G�0��K�yED
1,J*ܸ���d"܎&�G��Kh�d�c"3�����Bx��%����}w��g>����������Og���G��D�~I���E�浕�(b<�|�^z�����}I�:O�t�Ҙ�pi!B�x�DR��,�t+��5⑪zVE9]+�p��u��I$��~T�E@*�a�%�`ؒȷ�|\� ��Ϣ��|�6� �&@�t�f�E����PzL/s8��$g��w���y�I�Zs��W�.]�0�a ���!i}��ѥ�M�N���2���c^�(u�!"�l>˗;	��"�As�B$˸�j/0��;��5�	qi�V�;�!iUvwuG�EUQBU>'��B�qN6G��陖]8��k��?Z�-�(�N��%^�ҡ�>3rΣ�N<�IԎqc#b͖l�`|����5�f&	�6U2�.7u�}�����͗��q	�����`���>��V�gJ������z6*��S�Zҵe|>�H�f.�;U�n=v(
��3S�fk�XAՀ���U3�rCt�=Gk��+{F�>�"�>�yv��+-�6m4�ɚD�Vm�zZ����h���e`贅�U�z�h��T��!S4l �}oG8���Rw0{ͨ{֝3�a��:uܣg}��8;�B�>���q{�T�7�C���f`jU[0���#��H�N6< ����珇���{�tt�b6�;Jl���\#n;�y Ҡ��O���T��ϔ�-����6��]Ĺ�ް�א����{8�	��I��hk��6t%�l$��AƄ�d���
`��m���8ElXsᥗ_vʚ��_�=e)�`�do8����/
Z::�E��(l?߱�e�]Ɓ�?z{g��O:�ڃ��C�2�`��U�v>���7��o���(U��5}�+)�D[��&e	(��C��v�IN'���3��D8 ��3�R*β1�u<���y~�KB��@��*;�	�����L1P��y��I}�1<4�B�f۟o� B�lr
k��g\֣�P�w1�*���a}������+Z��R����H������Ё��'2v~��)����.���t�._n��{�?z�x�@�jSNE�-W.7��ԦWT�
0���jW�Ds�o~a�6	$�0Ƃ��!�I; !}"e���b�+��̥��j���S.�@J:�l��
�C$E�8j@�[����{���'ռ�J;>�	,ŋ�މ�Q�!�sY���gcGٚ������}N ��Τ�SJ�pt,PZ���]��t�w3�)b��XhD���V'����q^��r���?�W	8���Y��n�iK�00$��o|ߍ���8�g$�P,QI����IE‟�tN�/Lm�|�7�!�%y���R��F�B�ڵ��G9�b�յ�/Yf w�*��yq)E-hs��(U?~LFc'ً\�MJଃ����s���Y��E*��1`)�Jլ���9)Gc�OE,�A�
�z��Ɲu|��P��>����;K�&��<�H|�#���ٿRf���s�>����H���j��ڳ��/�cy���v�̼͛muu�2�dԫRo��>�*�jw��"���z�<W����l!,�_��Z(O�+�տ�/��W��'�0�Ϋ�΄2Q�2E����Ҽ��9��M�`%d��ۛ�����~9B� 5p�$�Ґ���W�8eF�,�}� �Z��!ƶ��^HW��18 �9��H�)�+]�d[X�T�vu��-5�z�;Jɺ��6,`ݲ�o�௅>��Ϛ��~�D���7�rKXc����VE-sUr9��K7]�����3�����u�t0��H�&6aj�����M�{c+>��+��BW#b���[yV�@��`��c���%���f-q����:��Ģ���rƃ"�PZ�gL��.�|8�D5Q�  ³xp�G�{�FC��Ɓ*r"�{v�)�̽c�	tML!���,_��
u�\�7�w�zˀ��+W�t�䩆����d$��gb��6�D�<#���w�q�S�5�󗽽��)f�<P@ø��DZi��]]fÇ�S�q������%��vvN���c2	��5�.\�Hj��p��P��-�bW�d��V�����G���X�E��|(�V�g�-,�Y5K0xr$l�I�GK���_PƁ��d���f}����t窉��QT:�=�z��C��(�hE�hD��lHU @�*��s�>�.�]0� �<�b���ޜ�
54 ��w9�%�F�#2�X\�=ڵ{��'5g���9��5�R5)N<�Z�d!ӢJ�&&�@�hS�~�3�Q��ۼZ ���߯k���?�6n�Ǣ&���/|Q��)��i�p��7C�������cȂ���S�.)-�*d�#�00$���WoA5�/���p�ctʫ�^0O��1�/4���h��c��=Ua\���s���׽��20�3�_�����!����)�O&zb�?�(<��7���-�s��� r/��3�M��� F3���x�6�;�z[k��3��"mtzxH�S�7����z�7��&mT�a�0��i�4�s�!������-��~SR��_R�.H~��^x��8�U|<�؃�"�
L�}����1	��	1
�W�B��d�A�VV��[�mnȠ\���oS���F�Ra�:yd�o�W 'Y��gu����=d�2��Ŏn���%7~��G���j����|���Ŋ��j�_GC�W=��3��o{x�wF��zS�Js�E�:��������B)���s��n�]<*"��k�Ot��Q�0�0�m�1��/���M
�3uU1�!��@v7E��(�bkؘ͙�xd�yCtݸ�����3���`s��U����%y�h�B�|������խl ���"�f#��R��`�F~�|��aي��V�6l����a���%�*T#�8a`��Z�2��p���s�='~�[����^ڱCj���� �3���s� ��A����;Gb+�v�����ꖫ�r�f���k�1��}�wD ��q�ݼRǼgA{�"t��,����- ,v�I�
c��|����Kd�yjm��x�����#�`�o��P��;�
=�[�k$8@%9�
��գ!�7�C\6��k���4ג2K�M䀣j_��6��d�-��F`��I���C#�g؈3�^TWoVBm��^ ����D?���'�9�SP+�ct��ePڼ�Y r>`{��/�J���@碲��ZY�9�C���V��2J(_>�ނ���]�fS��`�n��Ht;o��w� :WS�e�65&Bq�rg
5-Ζ(A pG	�Ĉy�y�X*�xI�ZEW
�N��m�1I�;Z�4h�����5٠����"�D�Do�n��Y3!J?�!!Ez٦M�x0RI�m�<���x��:� ;{'��I;±���- ,�ق�B �'859b�b����M��(�,����_�@C޼��5��LON	 0##��0��>̤��X����Kq��>��O�F�{�z�5��#zD����UVx� �`�<�����r�p-���]i\�֐'&��j횵��M!����@��N� r�阶�s�t��-�_�;��?$ׅEB��V§U�xr�}6�I������*Q�g�^-dvn�������mT�����͛�wYh׆�Za睰kB���ʣ�;���J���k�v暈���d���Q�X��3�s��uj��4��Ʋ�+_�=��� �o����<��_l��)���i�L'�V�g���)���+�ȫF��gT��ϥ��=�ۼ���Mar|Z�:��{*౱δ��wB ��4u��Z��[�[t�肝��z������D�s��>�}��m.�ՙ@�% 3x� �T ��X-V+kYs^az�^�"T��x]����0�T�Ι��Bj�ħ�K [ձٚ���d\��P����T�̘�S��z��Lހh�|��bG���b��j&RN�L�����3�{<�i=� ��W���y��ls�<r;R��@�W��IQФ��E!���lT�65�����YBֳAm�:p�hX��2��Bp��Pȉ
��%U�K^���>�p��|-��p�O����G��k��<�۹�,a�"�395��B�E�z��T}����~XK6��nM�x���U+@%�2>�  � �v�_t?�r�U���@��f-_�B{ξ��ú�:�U{;Z5�_y����0�J�c��%bFd�ē��Ƴo�"�Y4�(�:\зX�)6!�Ύ��p�%�]��ٙ��_�=�Ʒ�i����S�H/�������^{�U��~��O˾��?�D���>��e��K>�پ̾�̉�r8���p���:�(��Ü����yAiN:�;�߭[�F�ED�ݻ���i���U��rH:��C�5���������2����kr��#W_A$]�D��3�|��Ww���yg~�@/�xk>t����_ms�F�v�%z��OC��$C�\}��D۳<�<Y{���Y����Z�;Z&�ӳ��K�N�a@_�6� |���g�b���wd�Dҽ�)Z
������ �p�����B��j�>�� (A�j5ɮA�B|����TX�m���g~����R��
�Z��4��k�}�U�y�Fn����G Ǖc�l�I�G\{8S�*?��pah��9UhL������j���H��\�O`�f�0  V"�iSL�5�86tO����1����{����ºkm���J�t�9�V�L�C����R៞�h4����� ��Y�?���D��t<|�oh#��?=x�~-|6�ukׇ��Aa�Oi�����j����}��O���?��׾�����]?��t�F��Cw
���|n��,�4e���!9��űi/6Z���I�� u@ҳ�>%�r+�MT1�k$2�=�1���ѻ�R�E[&R��.�ba�������������,�a�ο�<qƋ��ƴꄢ�.!���%��&��3�yT+��"�ޣ��͟�;95^x�E��C����+��n���6M<��˖7��䢼PU���+�{��ɓ�c���e��d�����ArJ������3D��&���� #�zٖ
��K22|x3���5X�)�1��,Dn���ځ�7�5G��5�4��)��g�T�i�ZK{!F
5E���j�j9�1��a��Y[)�T��u@���s��4s,��ZV�W:Ί����b�lK�.Vf���S\a�H"�Љl\J��&\ϒ�'�hP�Tyۦ�f*���4b�u�Z�ٚ<5xJ�YΉc�R���Q�I��X�s�#�2ԥ(��Ŷ6���G%F4^4k,k���&���a�ɨ\`W��>z��K-��LMt*0�(�*}�{(� ��rm��a�.�%;}�H�>���-�thIڟ:ڔ��`���\6lX'��w��]�q�]�>��h;W^�E砨�^��6{�w�!@JS	R�7�ts�/���(P��7�LUۧ�;����q�i�嫐�^�m����N�BEZ�kir�CV��Ĉ�ج$���-ii #����}j{��y����z�ְu��#  ��{ @��cy�5�z�ʞ`'��|��m��,����� ��OL���Ne�Bd�w��E���c���M�]u!'�����������G��QP��c_����Z_�H�}���\l�GD�V��\c��kS�#�I�NU�'E���!��X�����= 2rzSС���G�f�q�O���*j��ߋ4��3$��.K������]�׼�\��/j�j/��<&mb��xK���v�����'Ak��i�S��ʃ�8g��˳4��$�p�Qn\���0ix��K�;��jT�'b%6P"w� �Z%����OuفQ1N�0���`sߵs���xZ���>1��a�!��"8}zT���;;d\R���-��Q�f�"o-���,~*F��&�C=� -Q�Ai����aG{x�	�C"{,�e�������2dn B���00Y������A��	L�/�X�3�n� ���5x^)u���"������ �Y�DG�7���F��o��|��h%BI���},l4��G?zP"� n�)xދ�#4����٫��kڼy��"�m�4b��[Z��L*ղ�y�xG��w�9 ���Jl�F����=m��=���*�ŋ�oٰ�oq����c�>����V>:0�a��U��$φy��J�׌�t,�>֌+p���Ew�����"�*䈽X�=)�ix�be�e�f9�&�hn@�����Z��_�<k3���S�0?�&e
lp��4�ۥ�Su�;q2�wny��Rٚ��@�Y�m���qS�(�x���  0�ϩ�s�4�KU��/��p(����{Z����\|�	�g����eE���А�����P�a�ٿ��)����rX���4�9;]�i523��t8ik����ȠQ�l!�\�-�����?�g��Y)�a9V��F���#��Q���WS���=���q˭7�f�u�T��H�� ���Kt�]���ZPa��Sk�s�yzU�m�'�� 
f���Ο
̈~=��3ᆛnל���k�O���!Q�x�W���p��;�S�Ы y��;�� )s9��6�(�� U�Jv����G ����	
Tbw&�N�������̸����}�~fTty�6
-:Go��s���������#���G��9�`��5j?�}�6e����5l<U˴�}�G弣�q���g�^��Ɓ��d�V����a���g_�Z��H{�\��	�vm��.����!E1�́�]ݽ�w&�fh�{�d������oY��졙�?��B0��Ji��X�M����9u�7a
lVCm���7lnJ��D�K3��ɖ�K*&��O��{[Og8�ʛ��s�`���`h��A&¾��
7�׳w+Ȝ	�^�lM�%�w/S	��kqMMO�A���S�㴈9r�n��Y�@ϔM�4(�zd���9����PԌc`t�>�<z�k#.�Z�ƈL��ڜ�ɍ7&��Ȑ�GB��XJ�P�Vlr�R �M牴�\cc���M���A/J隧�B�s���p_�-�:�V��-�{��@��C�=�ã�f0,n�,��o׍�cD��X�>^�>�����ß�ɟ(5�"�|g�F��D�hP����'	�Q���Ɛ���0q;�~@�����oڬIM���_����|���1��@ �5����%��h��Ŝ0E�f����J�k0�������W$�Md����0��lO���͗�+�
 ���8���[o����2�K�~�t� ��k7�7���.;+��K.�$�=��B3RO=����)�j����<��r�5 �CQ��0�]�Z�w���3�&�X�7Q��ğր�U��l���h�y���=[�S�]إE�x3����C������z̓��W{�G���˷�ϰ�B%��Yv"���9����_��s������N����=�;�Q����y;��y�m�e� T�(��n����Q�����g�o5�;�(q���,����|$�sg$�笁/H�Z���)!" �P?J�I����5�1x�H4��� R<SS���co���z��A�(Ld��щZ�!` Zȶ\��WT��o�p�=�T�$҅�u�M���&�]�J�PE*��K�)�}��7m}���5��cG������[Z���g3����G�.���������?}���C�ּ����K_��2D��`�c'Ȅ�=� ��s�M��L��= ��:�ŎN�ɜ�P�'-?��UG*s�������t�cv���8ƦV��:W���J�
f>�Cl3 ��q˭�(m���㱃�f۶�a������G�O���K�y?��S�M;{v:v���b�{�B|K�.k�
�H�qO�G~8`�(#�;qGNKbۋ��͗���R��D��[�����c��g��4���#:7QW8��=;�^:ȱ'��R��X%z����������^����Ii�M���}�0hϹ�n��th<DZm�B�&�G;]���&�|�m���Do�@W��A�7"e��%C��U+�zE�?����۔�8���z﫚]=���G�/h���SI'�Ă�jϲ>7+ݫi�`Cod�R�,rR�CC#���-޹�=��Ѕ�;:��紫�5�\M+�I��M7}@�XD�ؘ88��֙��#��ka�Qm���6yJ�J�X��5@�"0p�.Z"/��\.������Kڌz{�նoú��s�ޫ
%t��1�i�Nk#�?t��֫����5�R��C�#�-𺸿�x@"�\3�];w��^�'0���ǖ�PT>9���]!�����T�g4�Y���e�/���u�ݠ��5�l?���e0jwHD2���s$p8�ö� SpZḠ��`��QS��9��y�e��P���mr4�/\O@�y 
#�G�sc,�Ei��m�3�i:9���Q�V��ӓ���Y�����!���ͷ��.�=o	��z�89��({qS{�UƷbF�r�8�/[�s}�T���mAޭ6�H�h-�J��E��" '/�W�P����R�Y[���
G��8�-�� Ik�'bDs.ݑ��j��,��c>@<���MT%m=6�;*����E�~�વF��/s �(2w�1���2���jsQ]K5t���r�����@�h�2Ü�N3��3�	|y�@
���CI\:��̼�h�w���K�|X�n.m�3"���mH%�B�)e�Θ�Q�9�%���N����!Kc`.>��I}�8RJ^z�.�R������eO�C���ޏ?Zlm)�B��6O��C�UTDEPG&g@Ts,��Q�g��D���KSq����E����5`�6��<yL�U!�:.�`�گ2vD�(��ao�8��dϾ����U�*ªg�!�VK��K/jd��[*pt��A]�����Z6ftO�#��oW}|���/�>b�8����!=�X��?�nK���ɷ���o��B1��>���Z�Zlb�
�x>�����u��⹳�������vۭ�#)l>���:u-�	�Z�E�1��`��<l<�4���'�����%�{H1�C=b�[��jv������ۥxAgo�0���#�
͈9������ke����ָ2z���I�m6J�.�����u����L�g���[ uv�b�q
Zr_I*�9]�7(p�^IT{D���L��(�y0�����.��}Pb���@\������HUk�Z��^���=�S
���9jϥ͞_����g{mdO�"[Ȅs�z�_R)�Y�*������9〰o ��qp�ͩ"N��2�"+�It�]|��nM�!���y���'�@$)�<yM� �8��G@ʒA tL��.Y*� ��q��jZU�@G����]w�ҩGlB<���k޷o�@�*q$�i�Ox�����zN�HB�0�7�!z�����
���;�z��-�믿^��<9
M��D���s�Y���ɤ�\ �͸���[��B@�g��L�|��p&'����{��{�LH$c�h16DhY�r��O�*���-QI�1�w��Q��ߓ�7Ƅ�Nɫs�IrO=���sId��?}H�=c�b��j���%���θ�L�����sH�������ZIb40� �$��.���s 5���&��zq`�T<"p���y���tv����߻�����s��p ����?pȐ)D�J4���1$�|�,@���Y��( k��q�tƁ�(��<7�:it�>����;>xJ�[	<"9*P��hl��D�J֬����k�W?��;OO�,��K#�Q��{�zATcj2��+���2̙�7����ܘ�::�r
�eus)��i93&����@N!���#�CJ	�W��]c��f���%�U�_�_�\��׻�N*սЯ��02"lfY���H`@E��QnlьpF%&Qi�3�0����hXd�޲=�*:�#����KDQ��&�F*�������I��nE�W�u�`��M��j.��[У��Xl� �@�g�����b롱��m�1���C��u3���%b�zc��͗m�
���Q�*i�!�|�d(B��H ��.�ul��:�z��k�5����`�@�����f�!�	�A1� �_�ş���
p
EhӦͲ�85'��ͧ�4��'�D��)?{to�+� �d�+�~�V��?u[�v��_��@#@Ш.;��:r*q�����c%8��=���n�Ͻ>Ǿ�u�[�rn���ۼ]f{��m��N���_C�`8��k~�:D���3>�[�c� J=	�Φ9������ا���^3>:�v33���>&:�����Iw��{Y��ͳ;e�$p&��ۭY�t���番lL�p=�~�1�u�P8b����t���Ӯʓ���䰺
���YD�ȑ��]k�$#{�EER8�|-�]��������{�%'��:!� ���
%qD�,W<�9�]�(�I��:r]p2l�\i��7} �j]��Z]c��W6r%�S�>��ղRD�t�9@x��EҾ'O����v�t�U�F?P8&<l5�e"��SL�9E��ڴ��1	X�|g�sNƍ	F���c� �H�D!�XT����,"���?��N�1n�6�`��FE���'���x�ַ�ՐZ�J1j�S��.�M��zA��rI����x�Z���H�4eG�c������MRkV��0�3�i�@�i�~�覍�*<<B��3"�	���1� Q �r�V�ȣ�
�T������`�  ;w�y�a�c��@��XQy����"i�z�*�Q��Ǵ)��������i kl���qs�:���D�{`�(\���jsg���Cj�ĽPu�� C���!SQd}�Q��}S��BhD��5��gA�C�[X���7�ɡa�ߩj�X9qӲO�Y���|���#���K8';R;t�h��G���8��B=r��V���}a�=���){v�Xa��8��^�8��o'���IR2k|���翶���MEC�LH��V�* }AK�eG��ҁ+��r-���q6>'b�i?#�����m�j�3y� �(�p�������եZT�;�Q�zhPv �Wcd��vR�#��[�n������+�4�;���L�a�1���w�7�9�o X�� O��A�KH{-]�LN�`����ښĎ�ΠCY���ڧ���]c5?��p3Ǧ͛­����B"N������OnW�쮻~=\��Z�iY���^r�p�H[�Rf� m�`i��c8- Mv!ɋ!�e�����:�������A~&�����P���1��k|�w��3��pH]+�7���\�њ��C��k�U�v�=�(������י�`�!�`&u�!5�^�P5z�N�jd"�k׮8��b���D�x�rO2�<��K��jjrF��h�����������[�R���7�g�bM0&�����\K��8P�`ok8���/�l["����ꌾ�!�����=�C,ƃ��U-9U:�BY���������� �'���o�͚`,QU�	���C��hLra�oN�a�+����(�g;����t�45�� H$����K�a�I�f��ܖwabנ�ѵ*Be`�>���vIXk�ű���7&�*����gp  ex'�8�ۤ'FN�����	����w�t�3h����pp�-��h3�(B�B`A����̓�C��`1� ~�:J9״����� �b� �����}_a{
Y�{e[V ��D՟�f�������r�����F����3�M��(S�T�|Pixn�="��"sD�Jc^HA�:��C�����!R��F�'�04�ZР�
��|��wh����<5)���u�}�i�is��ĒתF��x��@�L�4�l\�|c��݊��Y�|V��e�>�`�i)d�>�!(2���
�c,H'o��j=�_���D�1���Bca�>5/�J������a<X�r,. J�zk���T�~.������̌��tO�*I��� w���ڃS�ZS�����FK+U;P�i|r�\�<=���	l6dg����y�I����Z�hf*9�Ȼl�����r֡�`Ϋ�6��k*D�Y�>�m?*�mn����M3�I5��@Y�]�;R7	����w^(�9��T�ͽ�	�,�t��HMX�S8�ί�Ϩ`6��.�	Yj����t8y��I�u�J3#]��]-b_*�H�*b�į�X#g2�m�q��hA���7�%0�����S�]�&c�I��i7���L�ϋ��T6Nʌ ��1C1*�S�>�:�Rp��#G��5�߰^�)��N?qH���g��n-�v�
[�\�v��=�th-<��׿xi������"ډ_��W�Rw����S	�`�яt����JK�*R��^�ߒ�v�%���d̒���K�ZJ"f�2٩HhѺ!��X���Qu�yJ{�]w}4�~�m�z i��|���,�A���5k��sE����6�����>�x�j�3'N�V� ��{�� �}�c��M;iz>�>��7����K���~���g m�����x-��(�BDz���о��M/��9q��1ʶ��<��I��Ie$ق����
h"��(SJ���g�}�g�&���vu�:FȞ93���9��}��ў#'BKO�2ϗ�7��@�Ӷ��gw�g�������t!�F��s�a8�&�0�֮���a��a���Z�����Q�֐0`�&=��Uc��ے�=i�	�����k5oOڌ��D:�Ѵ2,r ��L��͓���+҅��*!ݐĿI��0�ʶ�|�2mx�Lb@����e�=�{�:ĥ!}����h��t�G1T�ƣ
�+Ҧ|��`⊓���z<����{�+l��!�m��j|�������Dx�&��Om'��c�5����w��q]���=��[��D����-N&8���"�^6���۶Ka�E��W\��Z�����blH���C��4c�q| ��{��פ��&�����O*���RI2"!iËaA�;� ������N/����+b7<<)�1<��.��޳H �$>��c�#���Q���a�_d+xƧ��h�@:�+] �#˂Q��i���u8��U�w�����.��R�'��}�1�Ţ�g;{�\�����Wm�'M�"#�Y�P��ݖ\l�G�'�4����.R���z��B�=3
�0p����8��$�hͬ4��mLA��`W��Xh��;n�`��#�hI%D]�6�ٌ\6i������W��_]�ʚ���>5�O�W�c����]+��\�94_3�u���D[2�TL%VGgc�Ҧ��٣��0k�l�"�a���_��æo�9�����L�?���֌��Sc�����ϛʌ�k��L�鰸�^�����\�(٦@_Y*!KӡMݲ��1�(�t����6�2�Dp�K6泡ÀQ���jG��p_�g:q��
�C�a���D�s�`��W�O�c�z-n�y��Iԁɫ�9H���}�G�V��J��$����UE�jU�ڰR|i�I�eKW�?��y���u��~�]��6��3=+f�, V��	��E�T$*�D2�h�eJ�U��\�����C.��*�/�+NbQ�%9Z,9EǱhUHP�Hp�B`f�̂��޷۷��{��~}�g .��GN͠��oy��=�s�y�sl�Y������gԶ��[�ٳk�ȡ#��勗�͘=�BA@���a�Ξ?n���s�l=��¿��?�u?����:�'��1�Yi�qŖ������j�p�P�-~��b�&WP�'xP��Q� c�_�bx�� {-QT�,�����9��-�Ҹ��).�`�ٗ	j$��͑�Z�"~���d�xA����g�yV�����UZ�O�+��߯����v���r��h%۸��ٖ1�F�a������������;}��2Ec�ʮ=z�`ٻ#�>��3�ı���n�^�x)\�q����X��
��p~��쀟^�����:����p���,`94�ǟ�6��@���`W�!�C����74����6�N*�~#�+���C�^VC�����vf��%�P��wt�ʵв���sK�a�n�)3��������q�7+��4��\��\k��6�m
�d@;��7�%VB;��Q��F	��=�ʑa��a�|K ���"��^n�\ӷ�:Ѫ����]�vO����?'��\� �PKG3e�`V���Ic��}��'O�`�D���e���jSHݻg�t�Vl/�Rj�f���<ب_��{yy��� 3�9]��Q�s@4�#��Ճ1���(!���dYX�r��1�',c����'/�4��~�_����Yx����%���~*;zL�t&1�� ��|ܮأB8u����Z�L\�����pox�p2(�۹��xm�@81���T2?���)M��^ݿ��&�,'�vݣ:���[Ѩ���ͯ�E��^xA�A*�Jp��@���'M����EI��"M} +�g�:=�t�=a��@ݵ{����w7LA���hu���)	��� d�砸���@8��m7��!��Bp��eorm|�X�,r����X��.*��(� G�^�6K�J!򭈳�����׌`�1#�pUJ�\3���	�ɃӦ�h�K�I��r򲮃��<蚛~���1Y�':��h��T��" ҜT���r�<>3s�V��
'>� ڜd9��0��Y_��)�w��"w����q���p�6Ч��}7':u�͎�� S�t���U+�ꍰ��*�iç��{�+�)����21j�-�;<���o2�Vͻ�+��.$s Q�Vc��~�3އ]Y.cƑ
����];�~q6��)D~�-�����)d��J�E��-֗= @��Ã������4�G���}��K
���y��?��?Rt�'~�'<Ο?/� /](�a|R�3��G�L���������|�Ͽ"[�����n�|~�
Y�3����Q^��zƇߣ"�-��i.��:u���92N ���X��n[{.�_���I��9%�=b��Gd���/���E@o�9�*n(Fte��3fLwU�<�w�~3�F5�Ǟ=��u��lnNCI��g����ptD�"��Kl5�,���G�'��k�_�S�L��)mPs")�����j�Q4!0;�~�j�7h\r`�~����6�J�ω�n�μD�R�qd��8��,�}uhC깬�=�DD7�u��="�#��¢�/uN�Kj��;�ê����'�k�P��L�~�X�J�0X��s��8��?v ]ft�Uf/��B뀑���������M ��F�-N�XY��=U{�Z�nzU�t{بC�<�E�V㠯G#����Ʈ�����J�S�H���n$rϞ�jJ#Ý���}G��D�"��_$B���oĈm"��f"����P& �E@����`tU�+&'@Idk$JN��X�ھxj1��E`�6W��c��p-�[
?��?//�!�����GW�$@m��ê*�Joh�Kt�#�h��X���x����']- �x���I�8j��1Ɩ�h��#�Ex��}��B�,����>�w���|�5�잸R<x�&������D6���w����y�S�^W�Q��4	�NlS�y"�I��Cii��+ҜzwB�%���Me�iz��ق}��8nn⛧ޒ�LjlzjV-�T��TR,�0:h߭��m:�>˞U���ۖ�`}�������Ernp�A��m��-kzdQ$�����(�-nb�#^"s)Eq�bt��B��ԙ�a��$m	�A�!1�R? ,�(E���b~)-�C����4y7r*�`۹y�9�?Hڷ�N[� "����B�R��5���ю��x&ۘ�/�d��(���Qˬ﾿���5��O�
O�xXf�����5��X�ۤ�K�#���^��n]��?GZ�j�8���/۶mU',@��J#L�o��I���@qÞ��lS��P������+��O�v&
��1E�(��,U',�͂RD��ޑR�T��f��� x�H|��~<|��4[{Q��.]Se6`f�C��N�E�������Ķ��3�h)ZF��Cx�-�?���3|��oǾ�U��	��z����p���y�~��U�A:�?p�kɉ��%y�s����u�0ol9�&���/m߼���[l�(�>�6f�J�4"v�vC���X��֓Y"@����s�7 2�>{��˗uNl>U�D�����hx��u��W/�."e����9+8pA�s��F��y���d�W���k
��p�Ə�6�Wk����,��տy�d�Va��I��mU����-.�)�+� �]�rE{:m��P�x���/$�࿧�M/N'*���?�qa�?}�;�1ey=��m3���bpM#ʥ�c{�{F%��|+�m|f�p����j�~��)-�D?ţ��.mJh�G�L|��ٓ���<�����~rHSUc�n7���Duޘ��s��,ÁjYz[�rVU�;"�G"l���r��D��s�kL<�)�6C�p nl��X ���MӺL��,6����V*��t����Oo<���9QRՀ7RL|>Ǣ{������H�@��G����	)�m�%oUDZ��*�$��YP��1��ӟ�i�$��H��P6�� �g������H�-�����+I�<Q��I��1�ڻ��łO�~���!���d��� ���F�g��S�����T*�u1�2�Cl2�(�C��E�M*�q$z�yI�Xv'2��0J����a�	��c���vH�n�fe$x^	�Ҷ���3-Ði��pN�ؼ�u�V�v�R� R
Dp8��㆙*�-�sݏM��(�#��(>�l����/��6!�=�&�cm��M�4a7,قg�����W��A���mn-�("���9�7+~gs�����WCul(�����բXC ���dN�0�
��H�|w8�N*�a�������μ���ằGtϝ9�K]}�)M�E;���K/_�}�� +��߬�ž�=nW�rN>g4~-����O��潎��NQ�^�w?���H&;��X̂@y�S�7oڟ6�����l��b��C#�B�(EH$@ms�'��Z����QƷ���w��s�.:�9�Ǐ�^�*��Q�AJ�U��^�Պ�����(m���z�)55`m�c_�VZ\�oBjD�mU/;��}��"6��#�|����Bo����p���p��U�Sv��p�בv#�5\<�=��~�TG�8��]�צ�T�m�R� $*�nv����o��@�/��/�����[t�,R��8`�)dD���@��#Ղ/T�Ф_��~yʜ*��P����v_4S`�î򮐚2��f�i�~��I�,��3���jv`�P��I�'�f�s!�?	w��ӻ������_�6��zo{�"�8~���5��$�F�R3ӳ7����������Ɠ��鷴?2��=�d��Ё��k��So���D��_����$��
e�X�\j*kȵn�^1<�-y�T�{ְ��+"�;C�;�U"� [5R�x���F]�I�E^"����M棭n�Q#� }�u�68���޼t5L-,ݫk΍�T
�����M�8�H&G2�C�d{�-V4ᒥp���L����d�V?b��9!{{�c``DU��;H���5�q��b�k��S7�|K}-�B>���oɗtyLX׍k+��^��ع�+}�'ó}F4@��u"W ���=��K�B�l�^�ߎ酒�C��百;Ξy[�O�p���z	�p�-��dNd�$ۀ�&��j!$�BG���=�*��R��Tքg">���!H�x%r��4��ڀ�?��?�E~E���Ǟ��O�4����RM����t�}��-J�! U|P)��
����� �^#ڰȸ>��~�^5O���"
GA��xǈ�_z�[����u��r�����+ϑn.<�_�q��H����E �x��Ӟ���^A�g�2D~z�w��ҵ���c�3b��'�,�n��<�g��5<Z��R���9b�;ឍ��B�y!е� #NE���lBs@cQQ����`u@�c=�Ն䖪��CO@����M�&�e�� C��ŏ�����t���E/))��n7�L|�:$ܛ�汖iIe볉�U���`��ޡ�l�\�F��=Ab�!@����2��{��4�
���tk*t�eI����6�N2�q���<���5*�)� ���u���pd����@���vlKJ1����y�e�H��~��r�p]�Ps:� k���7�(ϣ>Y,@I��8�������Ģwr���5��X2>����2&}�A�^��	�fCk�:����δ�s��Td(~)�vVRg��m�{vn7���h��\��$ф�����
�ڝ�.��#O�n)��S+4~꽯c4D��J�"�� ɶ�ݓ�^.i��
�Uk�ݓ¼{���?��{H��3�_�uG�I{�=$G��m*��x����`BP�}��i��5QZ�g��Ǝ����v��AZ�]�M�D�N���Vu�!m��	*|���2�wF��cǎ��)S����Ԁ�_���"ܹ;%~<6l4�;E18��w��?�t!��~E�N���)Z�8Q�C����g���c�&Ƿ�ڙ}[M�}�-Ͼa�G�Z��η�?��}�O�)��%�ƻGݮ���p��[_R}mu+��G��+N�>�a�g{�M�&j��d�>*g�,#���z��ν�B$���Y�j"� X8�Ќ�s�l����Nl�^MĔ=H=�mΡR��K��Һ䝀O ��5TS��BEcEw"� ?î����v��)��b�f�P ����������������P2�E3�ʀ�8��������i�g�f̖��(6��Z�!	���;2���6de(v���F ��W��'�+ݮ�+0 �d背Ԇl�,*DJ[��*��m��jEQt�Hc)�����k+���DMM��4&�����ޠ	��6�הc�U|<�2{��I�&�c2֫�fѮ)�ڧT�*G;�B��J.�պWYKh׌�Ⴧ$z�D�����ZDΈ
�x�\�IȂ�Of������&U��H���R^)U~���e������9&�o��o��"�����ߓ�!_c p�\��"�MZ��Qb\۝%=#|��!�Fg��CHY�O�L*&u!�A�Sd<I]�j��*����Q8��������/��/�OŞ���T�*<���?�����<x�l��x���G@�E�7�Qk<{�3�q�����i �#��}���C�o��e�l:�_ �o�qJ�bԮ�{!� �"��A�z+3�r���C1��,-/j�a���r��дzJq]�ū>+��U�bו��\�ɣ*�y�.g���ю6�{5���[��!��;HB�<�$��)2�Қ�a`�(���8<c����VA�����U::smǌ(��ĕcW�^,��L� T2r�<Fu�u`��>�� �D�27��ܣ���c�1����V`��=��'��w���}����iܼ������I�F)�*	�^�߽��w~Ep{���a�����j�3�E<���'�ax#�w5DN�Z����=��Hۜ:p��<dk�.	����	��F�1\m���t?yv?E�/ӑoو�w/6��*��6`V"�.�}yq>�ha����O�a�^������yG�q��Id��O��T�1?���Fs8���+�R���*�._���5fku|b��[t���VU C-mm,+�ݱ��ƿ��YSG��v{��^��h~�cK7�ܾ��G��s��O�;���'t�:t�`���}\� ǩR[�c`:���k�N�\�I�?2u�I*$���x���}�y�]9��%����+C��:���g+���tye�ޝ�jO�����H����U#���x������T�,�ϰ��p��$�C �l�!�����Q��3N��û ��A�{O�/�B�^r�Tp��f#�j0�G �~�C��ǡ�Q@��9n{U<���Mԋ��C��n��4o����]���"ov$K�`c}{~1������є$h�q����5��WW6>��+�p_*R��:�g�����N�xţ?3��RQڧe /�)cT���W�%j�-�l����/�,��x��]zH6Q�Ӽҕ����i���SZ�c���:r�Px��?���D>S[<6b6Չ�[YK|"��C9;�H�6}�:��iG��f�/:k��Tܗ�f�5 �4~?OBї�����>x�#������/$��u%"����{�@�@H��=�� �����K�����5� �����4����AD@��l{+)<E �i	�"a�42����P�] �dL����(Z;6O���I�l~������T��G���җ�$�G��?�������;f�h��fqa�RW 'F�s3��(�C�C�h��=�V�|��<lXn���=��&("!T��I�f������R���*��S1V��n[�a�ΥT��H��R��[,/��i���7����0`0��?���*=-�c�W�O�qc�ĸ�W��b�"E�7�1F��\o�1XS��K�\.�ν���EM���`�[c���يt��&�x8�;�4ڪT��̆��ă�pgy,�K���.�� "��r��{��t�^�����=矶?(~6o,��N:�.9u���9�)Ŷ�H�,ItTA>+@s��M��^�w{�����w}�M�fk%�z�t�6X	�ca�\��Zw�SD�m~B����L����!lhfs�b��V[�|"���q]3{��9�_S�5<XQ4N)�>�aN�	x�񝧾��ߙ��%�@U�iV�
g�\*z��Գ��ǆ���?w�6�����Cq@�i;-ijnZQ��Q�B��4SS���437+�F�Y�I�\����$��5SD٪�3価�И��'�����ّ~���7�`���Q�.v�o�yZ�$� ��ʒC����i����'5О���7�(�:�uI�O����\������xbI�s� 4�PT�#S��"��zfJ�5*����z�E�������-�6g�^�tQ|�##��s-��c$�;�wy��9�OPd��Tc���R�8p(%��=@٭�����o��sz��y����4?[�qF�{m\�kMit�����ر^ ܌5`y�>7}���������|������+��W��@���h�r�!��J�r�N�Vl�Y+�I�Z�Q�=Q�D�f��4w��s�~Ukw��r��a"A"�J�ƻT0Q�@�g��Ά�=�H�y���v�@9��#��S� G�
���j��mh:tQx^T�L;��Zr"V��B7ET������B�]M�1�NxF�}��Q��\t~)kr�j�B��H*�cQ�A��1YL&�c.V��X����o�%I��I9v�C�<�ޔ���M�������bb#��@.?�7��� K��!CC�P �&��GM�I�:{&R�C�T�q���HZ��#-���M���'c����&)p�`�jr~G��!�����g�$n�	o�w���ա�u Jz�T�wϘz�o�g�Jiۈ�Bs��y�T�y�sB���/F��ZEύg[7�s����ݞ�Q�}�<w8��{��;��"eu�Q��Tu\��r: .�<)�h?�A�n4\����ݿ�t2?>?C�A�*z��{}`Ɲ U��
����^-�zݽ�Udz�ld�وF��p�ͷ�܂�����ͱ���`�8h]���j$��]@ЃS�y�����C^x��֪�ܬ	ҏ���-Х�go��Dc���)��쇥�w�� "�Yǫ���%d� ޛH��][5�f���+Z����n�:�$�\��{�������B�P��}�A������NP���mC�e�
���hK4�t��R���Ri+�?S�v�@��{Sa�9��:����d���L����3� &��ߌ��ԝp��	sN?��~_6�M[�}����լؓT���S�4��JblᨁfɢEj4��O�E�N$�>zD�����?�\�nφ�㤤ljQ���`K*^�]��V�#�}�b��0�ٟ��@!@����@F�= {Jf�3� �~�7S��=���s$�� ����M���ҡz���(��*�f�%���_�����+��#w`���α�k�Q���y�o��o5E�ޟ��_S���o��b
�މG�1ܱ}���H]�%�~w�]z'�q�� ��;rf��"$���^��oVe�W��5�p)�p�6�u="�Z']I�lE�Ҷ��
2پ���7�1e�X^ ;�&&�G�l5���1�P`>xPϯ�Ȯ��W���x��EP���C ��NAr�"���2<�h%L1����J;d5��8��UED��nU���R�����K���-ߠ�NZe�`�3��2ͳ�&=�y �qC�S��W��a�mԏ> ����}p�m���[�1�Ah�L��jR�Cꟻ��J��1�a�)�I/��)���Q���Ey�=�� ���{�hKAF]Z�6:y5�=݌�K�©�������g�� ����%Li�����q��҂"�'9.�lE��N8y�{���@��]���)�Q�� ���?�v~�kI��c��TA���]��d�ۄ��v ¨PM���+�����e���ҥ���['��-��M:�H�D	�2���ǋOj�h1�o��C�'�_�p�Yo{XP��?��(S0�vy�\���j����?�4>��������V�E��imN�ۣ�Sr��	��>dF�%�{���ӳ��iqk�+�ǹ3g����Ȁ�;Q�[;�(r�����0i�:u�f�;B@<��G��F"�Lq��;��Ѱo��_�P����H�2$�\[�T��~I)cP80zl��l�]�h���`s�T6 V��1������3��>���~/^���^�wM������Z`i3�x�f�%���&�^xp�DJA���3�N"�^h[FB�1�<f����o|��tz�VSJ�w��5��*����� 
eޒOiYw�zYV����_s���7��^�ae� ms�G����$u�������㑊������T��T3���-~�@�E�SAO����;_�x��L>����9�y�&Q�Jh�.����v�W��>[-y
�Kef�/pm"�Tأ������5����;�����Q��z��Nvs��m(���)�ۑ�[��vû�t�8T�fO��>����f�.*m��ھ}Rk89�P���O�nBS��5k�	�x�j�i�B���f��#��!Jz���02�E�V8dP`R_cmYJ�{��Z�6
�?	�Pdʞ;I�fd� 78�%֫9S�S��̉�O�{w��s�{��pp����3�xb�߀�=f��١�ů����Zh�&�>6=q)�C3���4G8?����W��X��b4�u������S�C��#h%�T�CEj���·���9���F$��-�s���C��i|�;�*G��#'��jK�Ҽk�H��q���{f�C[����0b�t*�	Ga��0fϸ\7po6�nA�0���۫�商 �G�;��unp�ٖ�#xf����#ˆ��ͺ���-��륨��4>���|�pP�������48}��7lv_�2�����r���2s�^��©�o�k6Gz6��"�&���n��f�v��ט.������&�<��E���dX6�j�s04^����ظM��p�*1+ec�+��#j�d� sJ�nz�  �ޤ./Y:���Z�xU�0���h�M�ݣ���I���5��������EO��[mx^3z3�Oޥ�Q�2-~�d`XD�r aR��i�� 	�iƧC�,BҨ�V�:����`sǛM2��7/p�e��uo��%�;���B��p<��(@ ��F��h��/�m��bh� �`|6��χɝ�*�"q1��~2�M���F�zD��2�<p� ���㏽/�m���������Qc���8yfx! 5�7������L��L=�; �T��Q���P�$�D�H3�}{v띐��K�`�ԗ�;��e����Z�K��[���1/��n ��8�SO�o�8�	�q�{�1��y7Ν\�Q�Sj9s�b���fi�f��=R�̸��P�S��p��Kղ��w���ڙ�Ϊ�b��("6��
2�%Y6g'ww�GV��TA�G��s����ag=�(����&��|���ݎ�@�+E�7"U]<��z_SN�9:�]<���\��|Ϲ��S�>B+R0�DN�RP ��7�2��Fm���~ס��w�F��F*�ϳ���LݭÚ��Ϥ�ʒ�8�(�ɼ�,
�4�tTrR�}��5���;�;2g���;4�5�����;�����cST���n��ܸzU�������Sc���k>�F���"4?���Y�³b�/����R�A�����)(B��bsY�iĵ��W�]۟��\Ѿ�� �a'�`��}ؤ��-�8�ػV*v�t.χE'N5�4��+����U�`�>8���_��?�����˰��h;��6�e��`�J'��-)�Y�)��oa��I���f���ۺU:�Iǒ����\�v�����A������A�'�)�8����Q"����� c<k�$ ݽ{���{��s��sQ3�U̯��_���qU M]�9 3��<���N4���`����\�G旫�j?e_�U����`���}|���:�.6*�Ĩ��y�q�s?�]�( e�%�Hs���y����+6���*��
wWTq��.'G;�u>f�$pG������(�w�������mH��QE1G�Q.��A)W�N���=kd;h}��� �U@xh�,४�(�b���r��t�x���6�E�#
[�1�$ȫo��͎���<;Pn�D#�I�2�Ga��Ç���,����^��k�y1��ݻv��$�F�{�x�������S��RR6� -�7^��2�  �ޟ���x���_��:��?�S�J�&i�� >�G��w����J�� O�W���O>!CA�5�E&�M��\��+=��"����(E��6�W^yY�û���	�� ��AV���'�|��X�z謁���0�n����3��9lcvTc��+�_���J�w���j�8��1E%\���t�ѣ���ajvJQUY��G�#��9��P�Xm�ǪJ���Xrn�	p���O��#�b)��m��I� NE ݾtC2�D��]
\fNP�HJY3���#�0����Y�R=��*�\�l}*B��5)�y�EEI���ڂIѽ�:�cv����9��f�y���%EӿaV��u�
E�z�:'S���A��+�Gķd��"b�ƍ�b�@J=��~�#ILU����:�?��AO�?*��F��l}̒=���/-���-��r�z����Jr��įf#ame�ƫ��`K1���b��N7��E)�4�T��x�-�/]��vn5L'ĳmc#��-�0�mQ�����\ �s����Sy!�k��1`3� O�|C�8�x l�?��-^��l�.���5�f���n���ZF���\�Ǿ=��aL�����<�c ��������@eD{�;G�9@Z;L�fRɉ��}����e� �$c��}�YQ�R�����X��y�s�5�����bsG#M,�59?�[�o*B�M�X��&Y8��jd���x�qE�;"�k������TV���������ٷTa/���?�}�@��˻���_���jA������G�H��ࡃ���tt�~�}�D�y4��c�TL8{2��p�N�7خ����ǘK~��1k�Kp.�+��qaIG�k�6�����u�[��J��<{㌠H=�rsT���{����|X�C�Ѷ��+���%���mԟ�^�Q�?�k��c{�������2F�n�af~9\�u7����	6\��{�$d�!m�Ń���⦸�;E��96�[�R�T�*]��6���L�ܫm�$1�L�O~�StAY]��RM`����뢗$�M$^���Ș1��po,�!���1Ҁ���@`-/-�����)� ���Y!.�Z�z؛�K����6+�eC�j��Ed����� =0��I
H�(^x���t�/�ˊ���`��ر��쫉j�\>�Y�cH�o�Bb� ;� �Ө�z6
dБ���s?�җ�^!3�����h����d� �Ϻ�)�,@��l,Ũ�Um��ɓ'��=l�N�`��X<e�,١��V��w��c�;w�:��Cq����w޹�M����!�����7"�\)	���+�X1����/=M[���xNށW��m��qs)En�FN��w-�	��,̻�I�,���X�^چ����Z��V¢�g'Q��y~^!�bӾ�=
(qsyc�9�O'�]��SZ7��<����3���L|d�y^���~-������.s���q���y�1 �w!r�V��*��H��e�ӳs_��='����q
_���_�p��������r����~x��4��=��^=�6'kDx�nm���P�Kq���'�ض�V� �ɉ�~a�Q͵�:�\�~|xX��� Խ��
�����{��ö��ߐ�O�:tY�zޮ�ӓ�a�g<�+.��Ixwp˱���akP��j�\�,��\_��U�E��k�a�{e��?Z1{Ŝ�.��F-�VS{\Nlr=$����'H��5G��*6K:�6Ndg��G���K����x�uq�/Х�(mo���z<���/�eA�"� Ź�ƾ��b�t��&�HE��Y�@%���E���_��y2<2$�'��Q���%x��0����I��;1�J�#�'@�h$N~���_��u��s>t$�h�O�K:Р#L�vt���n�!N����@D�Q�9��4W �=��n�G�q��1�d���9���D��g?'-h�9۽un.ŏI��X�Qh;/y�Y4�5!Vh7֐�	�/^wV���XQ{��I���w��xš��/��]�缯,�qd��
���&���M�#�j}��J8w�j8��^�Ť�D0N�����F�IC:�E�R�/����Q�F�rC���B���P�(`ܠ)J�N��>p���<O�:�T۪�ϙ=�����r���ۊ^0i	<L����v���.]�"�*�����n�u玴�Fb9|�[��]5o�m��T�<��:F��R�cP�J�D�������F ˶�+�Gd���lE�l��aQ�D{'<5r����`��r@�!j��㜯����pO����x�/[����sl���#NhgS����ޢpF�],�7dk�T1̯��j��(=?=z�t����\��^������熿�<f�����i�-�����_��+�j�m��M�MĎ�a��5��]�B#�H��M�S�{�-�<F�{����{JŻ ��s!��������j�ȇ>,9P^����4���r�8�8�@y���%�n��W'R:�)�<�u��Jk���rXj4�;7��ys|Z� �|ax�		��P��}�Su��=�����JC���@F@���e�NE�ܕP?TR�f[j�t]H�x�z}���?[��Eq�Z��L�E�;QğC�w�u�6�N����H|��Tz�/��џn�<n)׋:�~�8f�CiC�o�#��s� �_�� �}U����~�J'����=���]o�7P��59��C����2ZfG��. �M�;ȺTk1�ӓ�Z/_�<�Y(ٜ͢0�����v�-w��tgƀ`�ݺ7[�d�[k;@� \�����Bՙ��}��A*<,�d_�3���/��<�G����k
&��X�l��T8 �UW!�0P��q!�y��	}�����Yi�޸qK�$7�t��!`WdX�3bC�޽��j���ᘪ��w���N]�����Ú���ܽ�ؒS�y!#������o���o=][�J��$T�Ը�{�>r�G N��[x�E��rQ���6��{MM ���}Of���s�\څ�Y9�=${H�E��ciq���m��fJ^�{��m��D�����Շ�f,f��U��?0�x�M;q�}��׵��9*%��O��w)-Zs�<Ǵa�3�r�n���&�(f/ wcV�����;p$����+����ٟ�9�k�Gl��ԣr��q^��S)�Fj�8��<�
���&q���Nx���H�v�O�yE�]�uo��0L��������Ź��\��[J.����J�G���ɜ��ݍdb#Ûo_?�7}hGh�\(8��RE����klyt���N��U�C��+�d�D}�^\�{8 �:�&}Ir3Ñ֒7D$�H�S�o�T��"x'�_�pmX�H�p0����H`��D�����!�Ƚ09񘘜<��lO�e����l������L�eu)����$��Jy�lPd�����;��3�p�úf�۸97d1ʶp@+��f,�20 </ףB��m�I��&5��~H�������3�.�A&�x� 0��oJSs8=pdX���/�q���w�9�e�l���t?`A;~<:xH�pex�+f��t��}��#�p'Wc`��Qm8Z(&\�pE�d�R�v�^��{&}��rH6��� �@E��3���X�l�cꝹ���UP2�u�)t����D�QPH�����hغ� I�.V��Z�&ydSߏ�d�H*R� �Z��}-�5 ��N�%=7B�׷�pn����l�{������>�E�"��ZL��(�U�Q���z7�(ɬ�gQ������IZ�?���Y�G�*��	�e	���/r���|N�=�N�(�:O�G�+�"7T�2�/_�����q"�B��@2�z��:-��up�U-
�w�.'�K�Չ�tm����Ⳏ92�p���p�l���T�T4$[����G��q^l>���N�mP�9�ʯ��l{�T�-�)��h�ࣹ�����dlŁ�hMT���2l���� �c� �[�Z�𽱙CNò�<#�����'�TD���32-Z�kuϜd�.ϣ"9L��J�Z���<`{�ږڐ�<yJ�N& U��=l��=��Jf����G�l/�YQM21�E�0�\do�Η㸎FI��ERk�ط�Ѥ�S�g�Z�gQ� CJ�"�����l�2�A��Ν�������{	s�J1k� n��G������*�:�c?�c���O�)��{�}O{$E���EƘ6��R�+���Z\20�Zѵ�/d��N��gNV��v�@��2��H�`}i�U72�$#���SOj? ���kً�����˽5f
��;�BުpE��u-�7mϺ����a5 E)9�Y���f���o�O���IU�IP�	G���O�����z����h'm���7y�������k�>ۊ���,��K�f�o���C���v
�V*�Ў-���sΆW*���K��΄�J�������}.����E�R�]��$Qh^�{f��m+ �i��Hc��1,
 8х�hR��η�087��R�QG1I-��c,�wM�*�518j�t�N��Tû%�{ܼYi8�� ���pM�Y�\IG0�]�+�y�q� ����e���{\F��i �n�sT���`ǁ��|�RL����D�J��&�2�|��.F����z���0�eDպã���~�;z� g�#c �F���k��qnN](��ܓi�U�z�*G���'"���n��?�6~x��̋Eނ��o:MU���}"��󧬨 ���ClaՎϿ�����띮��Ɗ#}�i�%!�n[s�y0�S����e"�e�V+�(u�y 	��ߣf�.\�:�j��L'S�]ɪ��w)	aSۼBxo`�����|�ۇsD܎��F>h�R���b�������� �.�������f��$���L�ոQ�K��������Q��}���f�C ��^U������vMl�����V'ʉ�(�Ϲ��maI9�����`���#J9ޙ�
�D��^�~쩧����K�P[��)VT=VkCp.`�΃=�^���B��+���|�Eq�R�	o���epS1{<sd[�A�(���<Aմ���D$R0����e df T�7䀏}ziiA{���ɻe�;��ZȈ�?n�sQ��!��r�]����>k"��"��*�$�����S����r܃�g͎�$*u������iV<#6�ߥ� ��E6c��/�J�-̆s�>��8.{�0�M60�>Bש�aO����tF�F��`��N/.y֌L�;��-�9�dc�;�E���ț�����d� #��7��)y�<ƶmӶg޴}
�:�eT�a��k��V�[V�~�98g��$�1!罣��^��8��^l�)��u)^�tmM��R\�^��@Ư��Ԗ":O��v��4s�=��	>{�ֽ���3azٜ��Q���� ^J,����l ��n;rzj�PHH���ޫ���Z�u\ðT�Id��-���Z��+��fwmIz�)�'������r�4�*�u��T�����^���B�+�̢t�00>��ϋ�7�pb1J�pыLx� �/���%.���T V�p�6 ?�k�NY���9�U�74���H]�D�Np#�q�<M�qTA+y���B��y����o�"�O� �wJ�ѣ�S�>l%*��ʲ�=�(�-2)Q����F��jۑ KԋH]�D�6�|2�v�5����UO�1n�"D;>>�����˺O<\"�x�)U��	�s~�z9��z�H����@�H�aHdc˻c�8t�`��HSu��Db���7���Xl�@����e���4�q��{%u����?Ӿ����r��Vtp�6�$3��"L<E�%���a���^�zO�O��I�+"�R�D~^(R�!F�}���������b1�vQ�ί����x����������]�0u%!�K䔭���3��mD�
@6���A��ja:�s줕��XyG�"�+���>�@R.x��i��=�w�G[�$h6\/E�6EJ��0=�xf�Mc�G�����
�����N7oÛ]�EX3�j��Aƣ� �"�=Nj�s���P��r�u�h.�bsU��u�^z^O����;���Ka��GՒ�j�ޚK���y�r�-'q����}��[����a��?�lo�2���ݙp��+ab��<��A׭�o� ���;�ӛk=l��?��D�L��������^?-U>��Dg�� 9����}�;��Gl�CQ�����z�!�A	��=�a��doݺ��=��3�hTY�� :e�JC�6l����7�*�h�U��u�v0)P��
����[�����9�ԥ����T3"���,��9��It����p�v��ygiM���h�v��9�^�g�L�i*|��#�B}�a����b{��Ӟ�
t�"�ڜ=��u)���Y����s�0'������j���_U�h ��w/w��10<rXŒ�w�W��>�'8���S�9Иx��(+D��������n��uF``^��
�h_K�^�ѲZt�w�';O��`��R�>��w{��?j�:�-̼s7\���a��;%e~��O�,x0�m�����ռ����l�簤g�C+�uT�{ ���`,l��֍��F�V�Dn�0(h�(��zX��2�}i�WOJ��Mh�6<*�0,�� ��<^Y'���*W��O��q��=ԩa(�˃�*L)�Hۮ&�277��3�~�gU��/�У�
)��"}k�w9�iAfm��\ m��I!��h*���SǞ}���z�F����y{�6�����w4��o�����m�B��up  �srgO�+ҡ��ճ��%oR�VV$tM���Ҋ��G��ZT�1����L��T�)K=��n�d��S�y�Α�A���Ͻ�{ (�~���֭�Z��K���MN�=q�I{v�k4!��\��L^��aDI/���6�=ī��%		<w&;��؄@�g}5ܼv]EQ��l�4���=UKT���d��8{w�5�5'&mA�B&��}�f�o�Z/�o�B�B䉳�;
Q���uwzJ��?�?#'i�� "��Ã2Խ��J��JU�+�&)�am�ld�C���Zi�(�PE^^�-�53Tp�+��������7Ê�5{d�]6�������(��~����J ���U{H�m]e�KD3s���{���	$�O��sѐ
�H��}�H�8m𘻛"����&����-���9�"��\].�٣���.`���Qh>F@Z�y�=���90Ͳ��S����Xc>Pƞ��e)���5F܊K"�K)��c*��0���$!���Hk��M,	���:�*�vﯧ��L>8nܻN�=��¶�|4 Q��F� z��S��Xh�`����:�fg�ݵ�:?Fl}���iy��n��N��?�A�zmi�5iu�PXQ�`O /)`�b#���'� ���=*�0{�C�����a�`s%[ՊJb��=���t���=
D���W��O��yh����04:��4@�5<k Fy,�a���rU�6��̽�� �M��	s�[woߔ���U���[gޖsNtkppD�B�$���s�i�*޺{G�K����1/�[���Z�r�J��}�V����|��ѓ��g�a���C���8e�q>ܛ�g�:)��=f��Of�� ����ĸ�Q�5��پ}B� 3/��fW���p8���~\
�S�d�Ν?����'�zL ����i����7ƹ8��l��a��"����>K`@��6&������\��i�����Q1K`������B+����=��s֎2j���+uC��ݔ����>��g�����:����)R�}�(\ng~6ka��57��t����]�}��W�����&|{�:䅺�.;k=�zFj�Q����s�C�$JkHTd�u���(ɗ�-�Ӌ�1빨jW���%3���.B�hהBc��h^�0w}�.@ϖ��pX��@&fP���*�
"0/����%]�osڼ?�X?c��M3�v����M��d^\�q �W	� ,�vdRp=R�T�>��S� !�A�	�e�M�FI�a������Bǃ ���=�D�{��,T&,�\��M4	��7 I�p�y���A,^˵��U�p��M*;)�/͇�Mb8(���	%靨T���81���u'V�rx�qE�5�h��v������P�2`�g�������W����7P	o��'���
VpO4V��Ș"K����+�j�}zjNRE�7����䐢�p��'��G�ҕ˚DE��!��8��Ml�� b����RЃz�8)�����|�����6�w�x0�1E݉��%�%��4$�M��1Xf��� ��0�T�uښ�;�̰H�����7�ٷφN��ek4T�F�m���c�?�����s����ʪ�9U�"���R��8��˙h��n+UEo����]P��E���}���b԰߈(��S��[�&��3��;�n^��c�n����Y�����?��DP�g��� �O	І\�\�+���Vwc�s������es��ܾ�۟����ꢊ��)]�@��A�J�q�l?�����I�]��ڨ�Vx�6�Dk�i[�W�L�'�oKS�l=F!nwx�Xk��	p�Ķ�.�;R�ix��l?k���v|��ן/��/{q�jh��k�I{pXѦg?���YҞIՂqb٧lńZ��=Q���>|�P8o��6�.��������{QRN*�9(j��Ap��'3�4�x�l b�%}�,��D>���R�j̈�b��{����Ѳ1G-�U����^i[)쥥E�߈���6��a8,̯�U��L��ɹ���'F�A� �"u�}��Guͩ=S���3����w��=�+�PV*l$y�S'O�֒R�_��0Cj'�fTͶn��L��4ɓa��Y�`Ep�~�#CQIŻ�17pFp\T��gG��T�"'e�Ae����B�lV�	��4�R'���^����׻�:E&��N�[�z��r��s����4����ߩvl�m�vV��M�������Kj�y9�?��nG;�z���m2�+�/�;wV�,��W�y/���K�d�l��ɘ",Ɗ�.Q��0�\	���F���� �a��o5����v\U"vlq��f�=&�!C�y�T� W�ꪤ������PQ;��X��{ !t����}��)�v��G�`G�M���jb :S��� �$�d!u^.�?�����x$�Ù�c�o��*�Ás��;�W��R���c��$� 8#�|K܉���)��1�|�@�C@䏶��W�n��+E��:}8m���un�6�T� @^\[յBDP312&o�g_�G�����$���sB�x̤��Ó¨>��a5��
�L��p���;��x�-pM�#����f|0N���s
��8�׮��{e�8��pv������]������6hG�h�7pF�n߼E����Tx���k�����Ub�ǚ�?F�9���gd���<W�ś�{����I������4ɢ6`^*���u�+�<��:����+�KՒR#D��F����9O��͙�080��QnlL{�%]h��*�M�w;K�a�ӛ9r^���֣"����J�~�4�ϳ�"��x�9�)��r7#�S���u����3/���	 _$e�t��pw�"�����y�Z�XI���~_4��Әg�<Q��+��CM�&����P7��.K'�{Q������/U��B{����ِ�x�o���9Ȥ�pT(*�Re��9�D')\�,�D�o��[̉�w�Z[v��^޸uK�Y\X�n�
�����:�h�G�|fe���WR��R��K�-iN�	t��?��i῍Q��'Kr�W��ak�8C>:v���X�(@�չy�Nx�Ǖ��� Yd�]��l$E���:��$�%���΅{�O�ϰ�D�Ut�*�X�~�"�8�H�`���(�g���}�`���ʹ"�^��-�.�@��׊"�4� 3��V�T.����H��t�̽��AW���i;��"�����mFRЃM%�F��_S�8�����߸l�|-<�?l۾M�k�<2F�q~(듢L�2���+��+��ٺv͹�D~�_�Lٞ�^J�0�}s��n:to�2���<�lB��< �:=�q!�H���qe��BƋ`	Uһw�(�|�މ��?���^�	"�)�����>ԍ6�mz��8b[�T���0�� ���BhvK�nk�µ��Ώ��_0\7T�x�1��@��D+���PD񭓯�?�X`Х[H�^Jo]�6u�M��:��FT�c�Z�Ź�>1��С���O��Ҝ��5ۏ2�й�_ք��d�ҵ!WI=�u"�k��Vz�s�bu���R��?s
�����p !��g���n@���f�u��ᢹ}fE��Z���s�T4q �]�;��IЕ�]Ou@@��M��<��x1\k0V���I2��
P�Y��3��a��{�]�Z:0(���B"bn�-������:��I���1)/T�˹yEB%O4���Lr�I��ɜ� l4�!5߹sK�b��Tt�23 �Ի�����:7�kC�.KK�$�ʻG�g8�����;q��?^+i���Ӛ��W�K)U5J��o�7ϼ%m8E�cW��LLq�}��b����Gx��N�-�O�� �-���X҂��'?>����3L�h��D}M�sĝ6���7ʙ6B�@cm@j*��>ى����Th�7{Q����+��3��fm#��R7��_0^8q'���G;�X��_)���Z��X��	�{��z�:�@�%O]�}��^�ٻ�F��z�V㩤^��"�U�^b��&��D�8�&����p�trG�D׫tx�B�.�P�+"�U0�Ed��c�H���X�����, ����GS�+J󅒋�co�:F*gȮ�f�ֈ��C�J3�^�pE�U�Q�w�D+��c-�J�̎��Yc����R[<ݎ�Y���vO�E�ɤ�ff�9��6�m�����K!@�l³�Vew��E��*�����_�b�a�9�5"4�Vӡ�m�ճ�R�/2f�����wd�w�����L�g�{V6)U�
��Z�."uFƃ�
�3v����3f�I)��	�m�E�W�D9B6��Ν�r��-k�l�ۀf�����0���
�LxD�(X�������8~�� �ˑv�|�� {�F=H�k��Tl��u Ch)�T|�@��>��_��=̅�;���۷_{"igx�D�̑V���W�{{�aE�+��t�m� #Ș֠���b��T������a ڭ�ge��I]�1-����W&�O4r���]��Ǵy���n�c������?ߒFdu΄����K>E���Cg�S�&�3f(�	%��̦��x�;�P�1<w�r8u�rX�k���ך
d��{r��]e�A�As,�^A��?tU�` �a�����Dt��F*�^[7�;}OMŖ��%���暡��n�P�Ԙgus=4��R˼̶"��X�7��м줧z�Ԭ��=�LD'�Gۊ
WM�R)꾕6��x��IM��8qp�CZ�_�2D��<F'����ɝ�7�G�b&? �T���w�Qz�	��*������:y�l���Q�9�6r</�ʕ�i���ʱ�	(�!e�B��"�؛Tb�����Mu 	 �v��-]��d�gּ���J���P-�6�H����[:Y��W��Q�o��"��C��!�N/b���^{M���ș�%QIU���U�&Ubx �x�|�L_�3g�It���{�.��k�"g\�e}��yEKz������~3r��>�T,b�kM�D�����%[�D=+6;E��jE�+ɳp�;����{��6�`"������y�81�D�D������K��&�*��U�Y�-V�ID}�:��(�H\m:��~��k�,snꖱ�����^�|�G�ö��9u�d�gC%/�|�OwoӑT6|��X����Mz��;�+��n�G\�n���b<iU�f�Q��ri@��p��Vl�m��8�" �c�y��4v��{����679�A�d��0ٜ)Û��i,Κw�b��#�I痼��Y�_o�ޙ�k��:yS-�(zp��~�������HI��4��,���v��,�_��=����>O7��8� rK��D���j\[��y���Z��b�=����v��UDߕό��z�:(K0j�馢H��7�s.ɱ^4;�Q�:�uͦ]5G�����I��n�X�8T7�|�����3H#�}�FqnzV���������bD6��7������I�W@�s�+���N�yF)�._gX�o�|�Z�s�������\ڇ>�!s�g�=�"�@y�O8�K��0b )"����l�����car�v2qD�f��4j���Q� t���&��ހ���\���U�ﭺ��߱}i�(X�P�n{&�r�C����,�{���⨓b%�	��*��lu֔ID.�-�W�	O��	�b/-�U��d}iU��(���:�� ��M5.\� [�GO��8d<o߽n޾)�����]iԵ����U�`�xi.���2<��ϫ@R}�(�R�TuY�g#�u|�Ə����Uހ�h{��xZ�9�v+r���s˾n,l,Ůs�@bEN]��ZTV��|Ѐ��io`8L�{��sf�G̩e2}��ۦ�jPV&�����_eЅݛ����o���_�r�M8�������:齐d��-h��r����Sx����w|D���B��6N�oG1\-������ݍ O268�Fb��z%vAI#�Kq�cuO��i�R�W&��?���K����4%��ۋ*ؼ��Hi�̯�S��sn#Y�1���4;T _������l��#[�u��`r���	<��;��*�	`�[yj��J�1 ��7O�9Rċ�Y6�ը�G���]2��FXDjw����!��`H�rh� �3�SҸ���9�{N����b��P�*�XO2uhx#��<��c�5-IRA���]�j@���H��H�����cq#{p/�gX���w1�9��r���]vÉ�J�<``�u�w_@HU�&��G;�dJ��,YlA�K	�u�4N�# w��r7r7�$"t�w�Dlț��bKB���+��R�a*�鬷���V�k�f�ͬ��3��@��B�EK��S�y�x�j��W_Ի��c���04�+䵒wLI�8E��T��1��~/��<�?2g,����]�*�� !�Z\�x��=sQU�Y��;� �l�����_�?�ۍ���+e�?�RwK�T���z����al���7��AE����b~n�3޹z%��7���Cel��a�6St[C�E��o�/ͼ7�]�Y+~�.2>:�����W4fnO7�RTް�#���mV���N߶uv��>��d��Q��h�ٍu��N�Ԗk|�\]2��-\7ص5�M��r�J@ҭ��p����~�a��tC�msw��������D����ߛ������6��O<����JaBsA��ڵ+&8�H��ؾS���{��*DI_c{ GΣo�7�8�6�Iŗ|����������J8u�MEВ�-:��;)2�7#��M`�Nf"y���Pөi���JlS����M,Z��Mo�cǏ���=TS����S��A z�2v�C����h�������;'������o��p(O�����m��zOT�9L��Q��7;z���T��ϋ���o��M"���	t� �bǪ��D|��*��N�Vd��0���_K�&�cP�F��lz��v[�p�(��H:g�;�1Wؗ�/Pk�R��U	�G��4�Ō���4�3 +e�xό��Pw=�R��,_�I�I�DAZUw������g�Uzo��f�Q�H�籸.d}���=�,�7�g���ia3*�S��F����[�P��� ��G�>f�_;{Ҽ�w¾�~�{%��X��1E�(e׷�r�:���zz�2f=�zd�Rm6X/���4t[�)����L��"�I]eb%�A�P����?���2�� ��B)bQ3�H���r]~���2Wj��z����,�\���@�O$rx<{vN���R�E��}X�N}qY<�j�f�0Y�)!�&��[7$W�z{�y�䯼�=-�r%Sk)�� :��H{o�6�	��ٷ1rh���N 9E�Gr�H�:�3:�t	���vf��p?��5���W��n�g���w_y�p�TTb�mQ���&)k<{ �3�p��1���2�+��Ҋ�7���R{:�#��:��,ܐi����
�:�9�;߰>��O�����7X�X'��X��o� ^$i<�}V%�8`�Jt�,>�<=��Pڤ\n�ʾB$���c��8�'�U�y������\�J)�J�pb�/K�k�l��"S�G���l��E��� J���N<螺?�s��\�\eR��m�j%O�J�<��/������>�Dl�8$[�M��5sΩ;Ƒ�׫(j��k�@�;[[��l�~�s����S!k��r�-ՈA�8섏<v4�w����Z��7l= uB1�(��a.Ļ�.ԋ�����K�p���V�q�����1/��R$'���YX��r��զ�)l;ǰ�Ņ�9EVx$
c8�D��}̕z������K��ٛYsJ�����iw:f稇󗮊W>^7�����VVՠa���H��bsu��Z��X���~�گ�Z����	gΝ�>@1���#�
8�7�]�V~���Ə��ի�b�A]�����`?v}F돔�<`�HA��K��iH�ϼ��R�-��d]�xYNo�����6�]ꀃ�>��V[dH�������B&�M����ђ��s:�_@N��j)Lػ`πW�8� y�j��-�u�jy \�rM���񭲕���UU�r݃��[
<���ҷ�%�%��	u�}�����e� �m?P�zC?[��ST���o9�޽W��2op���߫�
��A�� x������s�9;dᖖ����=���<"���^�Z�9A��l�f"U ~'��DM��^'������ɟK
%��UvG�-�Ht/y)��d��t���F��k�.��sݶ=�S�
fͰF�)ת��.N����1,EF)�4��Ijj��I��r �eX�>�eim%_���{𽔋���\�rz'X�jɄ�($qz��"��
�J|`Eu\i�ZU�-��oq��>��\a�L�`�c�E�z�8�Ő��şDl^\�::��7~�7�1��� 5Z���m�l��XyɎ����-����h��&�)�eE�FU!v�@"�{dl̨%���D8�*`����Yh{��ѹ�����*�H���x��CB�9 �Ώq�u&4�Rxj�52�ߏ�ޝ���"�K�5}|t�f.�sތ�%5V�Z�D���� M��*w�YN<�|�#b:\{�<H ���ƻ��(���q����7�Q=��:�g΋�`c����6@�އ����i�^hy����o}W��9����c�j�o`qs-��� �l�y��1�.;�F�^��I;�>��������W�!?�6OKEjz��#�A�~X�n����<y�"��h���{d��m�ڥ/2ƛ�j۞�w1@l-����z��Ͻ|��0n�<���X�a���0��jTEi�<Bَ��0U�f�� �����	����j*�HT`7U�B}uM��#�L '/��vU�\�]_r}:8�:Km�� z�!��b�2�u�ʝ���m��{�)�lsxߡ��~����M�$����?�̈�}��k�z��7��`!˶$l!�ц� #l�4����3^��a��<��`?��6a� �ԒZRk�M]U]��ffef���rc��;�DfUw���Χr��q�������{�=x�>�/ͪ!�;�=*J�m�vnW���gs�k���_���1�!W��3Y�S��C�+��lJ���SSK>�c��"�7Fr��zU�]��3�!c�[c'����B�]�Y���O۟��!�@C�T.��JR�J�g99<���2JT��D*M���2k�������~^)H|䩙E����{m�ڣ�~o��e]�NwS�ōf.�7��X06+��#eC�������������3bŸ�m6��1Q�jO5�t��~&�RȜ
��fx���d_��>tXv@J� JZ֢������b�O���Ϲ��o���6`j��	:�eg|}�Ǝ�^�����wK\ ��8A	�R�r��۶(H@dNu���I����26����_�2�t6��)�W$��'�	|����=��c��K�<sZ׋3�,v����GQ�Ų8fs�kV4Fd��m��.;v옏��MNLi_#"
��v�+���E�FZξGM��,댢}�y`x4�N"9��	%VI-��֒�ϟ���N	A���'��� jM�����bM���ˇ>�A{�;ߩ����w�
�F�p���u���k��/�6�X���fS�P]���W�Nڹ�+nu�X
M��@���D^��-D1��ǔ���S�7���ӟ�p�LH���@��D�O��_ܠ�hw�Z���2T�G����Щ�����Z���f��s]y����G�4)��j�� �^f�udR�ʥ���)�b����v�%�MW��.I��MǨ/�{����/ٯ���G^�J�^�ԙ�g��
��*�ē�I�W�G �d�PBw06ݰ��E�}�}�R�\,ۤ{2c[lp&�=U���k�<s�<F�
,.  )@�ҙ>����ٕ���PZ"�o3�"_\R��j}I����.8�<���(�j5 �����}�m񅂇�����	e6�G�k\��Ul���s�RX ~��.Vc��O����un�����I����J���>��26���oׂ���%E��bg����Ј��lN�8C~m�]p0���V�(�A#���� �B����y�]�茆.����������{��rYs ����?��'
%��	��J�q.�q�E�$����M�X�{2Hj�8�1�<��u�^�c���8Я#=�pъ��t�i�]�����V۶��>G�h��=�n�{�=���MF8��Qi�����fzD�A��2,�xm>�7��u]�|�<��r'����ta�^0k�����:c3�d	e���uҍ��ʬ���b��L6bmaɁDE�%bG�k���7dA�|^�|�׳�&�b�wsI��b�L&#N�r��+o~�ܱ��_�1�����W��]�_\�[Ʒ��yx�υ^{۟���i�3�{J�\[&0�΅f��#��5&v���k
5���E5߉�7l��܆V4o
���<T�JVI�; t&��@7¼��:���kց���o|���ߵ��n�ͩE�F�Z|Z�Me:r�P���D6/��|G-l�Yohp�5@����?y�j>���#6�_�;�h�h��l��2�t�9�j>̫q&4���S<�42�4���{Y����>i���N;%��3�7)�M3F���}��q�fA6��G��w�}�@ͷ��-�M׶n�m�fx6QR��'h_������{ﳉ�+�F]<�mͲ-ۊ�Ƨ�����&.���kR�al��vea8t>}H��h�&^����966�Z}�Vݶ�,����ԛ�R�52wH0�:uF�Ajy�U���
>���C�^V4ud|�n��6e�nٳ�nuǝ���̓�cW��,�N�k�Q�ʌ��������tt�8q���Y�>>�  �ne ��M*A��C�8_������дHcǲ>�>�B�eY��wvzBfz�v&����:�}�`���2=d�
lQ�Iy�[�����s� �~�~
]`s=����7 �pPC��3Qr
�+��:��j�K�з��m�s�)w���M��s�-�;l�B�:�w��p>���Y7M#C��Y�d3RcM�l�1_�םڿ~�C=T9P��ps7��IE"F Rי�rȌK�{n��h���F�����q~g؜(�o�&.NCR2�[�:
.����.EI�O���h~��S}Y��5v���Q�Uyx6��EƖx3��G>b�>j_��C�_Gq�P;eNd�_�Q���\� 	�SGAMK����k�Ss�a�Jm�T�S��j�哱�I�4$Y�D� ���#�&��H�������n`���\G�R�C���#I]��<K�g��'���5;� V~u�����sg��V��&����`P���N.�D�i"�� ���s�S���"v���,6j4�,4"��� ]d�#��9N?!�~��6�G6x�H��pb1�U7:#��G���AE/Kn�=d�n����N��}��PϦѴ)7ФD����#.���� ��?��'o��H5�82Jg��d.p�-��#��$�ځ�-:>�/�S����z�LDW0�e���ŀ�ns 2�%�E��Ҫ}��m֍Ѡ��~�[�<֐�j�����י�F����<Bw`
�E���S�aZ_��"��:]	*�ͼ�s�\�%���Ț�2�"��7�J)/G�tۚ��&���>�=�D\�w���{��`��"���͹�-d���4����d*S�j۟Eŝ��ʢ�_�jՇ��8��w��W���u�9�K6����M��g�u�e�����K�|����f+��l�-�A���H`1ECu��>
4f7�1&�;A��o>W#\m�NH;']�u܁Ѵg@�`Dw�:Uj�|k��7���&��/��b�FR�7��u�>:n&�is$2G��]c��l���r���z|��WK�H�a���������x�j��ſ���=.�a���"�!ڿ��`�4j��v�M#h�urvuX��a�ĺ1��i��c����c�5���bG7٬���+˫�������1Ge�A�ի���ܐ��z [���3vY*#�m�i��/�>3w}A�
���J�2����v��Cr�a���ņ�u®�ܱCY#�?�!��AEx� ���P�նs��թ���eN�:+@�w�>u� ����y�@)!�ܲSd����!��������xp}lه��d����M�(2s�[�k4b�_1֯6�g�N�2N�W,;��Aţ�u������x��I 8�<)lJP�ZZ�B�-o�_��_�R9�Y�F��,�ս��;�k��X�Q��BBq-`)Թ�f�������4��5�f22�9�R}VzD(�i���61��j�o>�>xO"�$�;.-�on���ꊆ�����Cv��򗂚��$6ץ xqz�V݋�28l�s��#� ��DP�d-E�r	�wP�uϿ���Y��H�y��4��RP���\Y�U247Ӧ���>h-._�|�ZL2B�)T�@��(�|�7d�sm4�4#�2�)	>��T�82��P|����Z�+��`�b��ZO`H7IE�#�ZxL�T_�768S��!}dC"\���iy�x΀:���r��s'���hj�N3�.
��` �7!z<�I�s׻\�ℌ��ۆ�=�OJ$Y�H@��z�q˱@}||�N8x=}��@�H�1Oy&�Ԩ�Lw+(�8=}ݞy�nJ���yr*hw3�;}�S&0��.�$�^���3�O��d�m��V����;��}��ѰN��(��JAV,�^��EMb��u�=���Q�I�d1!Ś�>yފh�ɜhy.\�l���	C�S�����o'.Y��%5��de7������Q��Kj���-"olT)�(v	��Q7E�6�ǆˆ�M8!�ӉO�0�G���%5�/~�9�z
>W�[��V~�A����z���e[�z���+o��ܙi��\X���+���s9�_s𲮆�2ҍ"��4�m�r3x��%[��{{���5�����;z�7%�y�7Y+\��S��;���~���T(�H��o30|U�O�cHG��5_�SI�����(˖�M�;�X�����q��1���jF�Y-��,*���ݹ�@C�ԓ�Zq�A��F�>Ⱦʊ�*�
n����}{�ۃ��!v
m=�kd.M��h�v+@����121	D���F���rt%49G��2rv��E��w�G�@���������I�b�����PQGsE�:���U#Ҵ����|�
}���+4�����a���~���w�W};Q�~H :�*#LC8^��li`��Fk�����y�ݾ�Y����uT(��)����w헳,*68�VWTz5�`�v��9_8͉�+LǶ���4�_<<k�\V�p�5{+�}��:D�do�dR��|s��mv溝?w)4���ڹsLҶ�ͥ@�����*�?9�6X��Q�x��%��O*����m�$�\(���q�!�t<z<7�z�$�@p�����%k���%"s�d`�زu���C>l���~� (j���Ϙ����uÜr��8��E��@V/YS��YsU�9�[��|���=rx[�Gn�|��#��X�V�"lNJV+���(��I����&���b�20|������66w���qk��Y�^��&��Y'z���в�0��/�o��ٳ*N&m�˭$��HuH���R˪�l����8��AJ\���S��fqp�T�#�N@KC�T'mޠU��R�v�&��(���}�~��~-��уؙt)�g�O��>1�N�R�Fd���OJ4 '�xŏ�����(J��o�C��s 3��rHE�Lʤ�B�.�"��G mpMq��N b��51n����c�v����n�~eQT3�3�%�$q�V+4���6/n�|�V;p�����!-�J�R�y"�����}<y-��? ����Y ��C�^�޸������cn�a7�"�T^�����,c?*ŝ��I��4�3�8\C� b�1v<�)�,��-��f5��|��ש�4���>D�6TF�g��@s��I*��_���N�d�$��"��=F;HJfn��n��993k_~�k���_��$57�g/ٱW��w���X�;k>v���$�Z�\w��]t�G �ՖB��=�M8p3��^�\�^��H�ϗP����M��!o{�6J]��+�f���O�����&�3�c��ص7�Y���}�+v���?�Ə*���bH���X/��i�D���
� E�0:����n;�Xm�i?���a3�p���7B���)R��)ٱ\�BϵsA��������n�t'�sPoZ����M�ϸ�:��a�*t��r�W��N.2T�}��!�9>do<��A��[�R�>)D4e����&��j����a>b�Q�"�����%ߠJV�����z�Ҥ��v�ݺe�o�����?�N��y�5ޤ8t�9��}�f$��5 g��%�X�6��F9�M7��q����`/����=�w�}�<���ǧN���'��R��Q�����U�!��y�G�;��!�Z(�"�E4���5�Ec��`W&'&��� �\_/@�G����v���j�U|�c� P���CG�ŗ^r�<(I���z�� ���6�F�{��瞻��?�s5`��_������S��}Sox���8��)H���o��,-���pRA���O�L������u�/��Y'#:�R�	�`�8��� a��x��G�9�c����(לx�y�	,'�� J�ql�t劽��'���G�(hy;0�F�&����b8O[�S�rF6�����rQ=��-����f 1G��O˳/�l�~���b����g�ʅ,�4d��j��Ї^���v�!Ke�7ť��Ϝ9y���F�����\>V����Bd��@(*M֊�`��R��Y	������u��s/��/��a�_�0HF��V(�l���@��l0��2I�/ 
v�		+}�d�T�1�FcU!zjԅ� Gb�,����:g��]y;Qظ� AL�4��|�����~U=&1u�t���#4@����I��L,�/R�� ���,@���|l�	��D�R�� �('b�D��HE�x-���e;���O�=�����a���{*��h��N�:BY�У�<�L������Z�k�a�ՆA<{&D5��dn<��s�ۊ��q��cy�av�����
���:��$�n��EbJ�����\��8=��z��	P����*KF75�����
��ϙ��r�Ԅ�# �R�\�jKtjBI�c=<:"G����G��Vd��.Z�T�E60 )����?�v����s�CM$�=�jF/X�(� ��v�!.�B�����$�|���f�B�2���tQ��|?d��gxt�Up|���m��Z����y���hR�P�ݠS��W�(m�G.���v�k��{C��_(���q��F=�JV�a�\誋2�����C��w�:����b?��7Z�����!�"�$�ymƟ�{�DA ^^\^��*��#�#�x�>�O��}��ߴ[��n�}㥡��sʣ;��9ț�5��
��Y����3q��B8�99:n{ЗΉ˒�L�k<v�	���,I]�<�N���^VD䡳���J2n4Н4~)���׏�mn$K��葃ۈ��(�ۻ�؈@nz��Q></�tk��9�u�h��>��s���=����;Ɔ4�t/K����H�E��<(:�Ъ	�K�uM��Ã5�}	s�mɹ�Y{��i�2����#6�4/#�ݜ���K�4_R�y5�Ĺ�.5���r�	�~���������xG�Gm�ڤ�2�����m9 �?��?u�6o��GvE:z��[]e�P�y�=����{��D+�v�}f2ǎ�v4?�'���r�z�:hc�<2}��O]���n���,�
�7�2(��m��!��|x�A+�"�W�)=��B.� �$(�C@�jϞ]�쇔/!�p��Y��W�&��f�-���8l��'�@Ƙ�ow����"�#G�	��7�&��`�P8)�z}��>��#���}~��!���'��<�e$�Z���Z�u�C�?&lme�2��S���Ґ�=<�7�b�
�&�r-�
�d����ao��W� ���:�=A�B!�hbYS(�Kk[{M51���v�T(��Ħc$wH�)��7�bS˫�Z�%��BEb!����A-8�I�G\"q�S�]��Q��N�F��.��)�ߠ���,��-�~(
7�\��Յ.B[��[r�Y�뵡^p��Ԙ�ڏ�U7���ťu�B�L�,<��"�<8�;��,�L��N������V!��D�M�[;���x-Q��� #�v>#��H�҉�ѫ���_���\�+W���P�!(�yhL�E�����WV� �>�J-L�um�2�wa�.]�\ґ�M ��fG���Cz��i)}��=�T�Q3���A �������� ?� Ɍ7�?��kÈ����pW����d}}J���a��#�;-�FcY��h(15�L��Ƅ{�[��6�_4�.>�7��Ly�Q�h�������{��]\���(��x0� pE<�~�Y�8ӔS*��>t��Jhv�	"��L��C���sW��"��V��y�l�G�4�PR`�����]{��ߣu����M���ڳxs*�`��zT��
,DRw��WVd�ǀ����A$q���P�`���=%-E�L��W��k�_���A��'�����}a�_G��N�[�ԇl�7]���oB��sH.h�ސ%,!����%D;��%�EJ��;�M(6fl�>ge����c����7Ч��>$8��Ȑ���l��!����Q��9}Ic٩V����-jw�^E�[r���sWl�NFȁ��͕{1~k�f�K��b�/>o���:K�Lw�g�V���X[�q���5����̵L���"��m(a��:�h�R��̀2��;���*Q(�9(�L�\;�	�t	�����Z5�e3�CU�W��x˿|`�4F4������ߛ4C��;�I9%�pƣR-Yi1��ĺ�f���*69�b'�O؁;��y�~]ΔlIKY$��FZ}�q3�f/�!Q���T�:�,�B��;�����g?�|9���Je�8x�vcߖ�C������EF�i2��#�/�.j�9 �*2:�:�һ~��Z�Ug�H�XS�G>_ҞB�^�Z��wb���IQfTc��x�Gvw9R�!㞈$B_�JS�I�ݲ]��|>���۪�jU5��a��ȷ�;*�F�cR���|��Vƚ�1b\����k��
�=s��]�17����1�4����~�R�R�Y���9��({�)ef2k��9y���E'b �-�u��;{W��L��>��k�zH,ח�� 	�f���A$�sI�A�.�E�M)p��@.u9�B�������VN������;Ͻt���h�+�/"`QT]b�&��Գ�!Z�a���91�W���V?5�)¹)�pC,�ΟB$[�^�PҴ�Nכk>��'�(EEr!���rn�W�ӌ5Z�8;�`;�G��ط7�ro��[$0�� s"����DY����@'��SG!-(G�r��.�P�����\ȇn<�<�� 5�����;��Ï<�@���/��/�4�z��� !45��]��&55��O�����}r��kX  _�/��ȧ䀚u<5��x�����-��U�!(/ y�� L��Rڛplta"/5X��v���!F�(p�Ls�E)��(�^P����Xbh ׽�=��߲(|0~xG�ѡ�C���� �����T&��1�/�K_@|���gC]�?{��pP���<�s�ý\���-Ӹ�8}&p[�����`��q�3�ҭ�9���߫���B��P���>�7����bf�3�t���������Ej<B�`��-��6�B��	̿���t���T�N�g5�	�2@�/)���t�&g�[�z�Z#��k����Uq���Q�J�RV��#ie�|��.Y#ފG�t�O��Y�%l\��͍/������cL$�'PX�nh��P��*����s/���5�9���c�<`���)��Y��T�v�҂m�2f�o�������xm��mj�K��=�������F��e̵&��MO�"�����¶�ܞ�p��}N�Wj���y�R��P���6�ě���&O�v=+�W����H,�ZC(��[�9�#i������f�1�
�E7���;]�}s#�F�Y6T�-��'s�@�#b�v l��Ɇ�����ta��P��[��;;j���0�_��"D����,�i��p�:W��U���r������Z��$�aզ�����K68<`w�6�k?�u��	n(lȽ�?s(���#Ќ߱c�}���������S�o��%�Dc
i��k�oo�-#����% !�ml���8�ox�ڛ ��������4�@o�B#�>w9v��A��>���<\�R��۷/~[�Q�/��g��]j���64`�ᛅ<��;���!���/�f~� �v��/46��,������x��)�M���F�b������g�ͬ��uw����6����=��v��y�:g����dmL_���+���БW�踰��j89S�7،�Y��۪�('�>91�(��y�"�ո�:~!S�ds���uF�+��O}���w��S'�7'�H�yN`4�E�]D4&L�r�b����ȗ۫�uw���*9j{��\��?��;�=V�ju�v���f�C���e(m��?�Zo�J�����'��STI�=�FY��u�8n ��؝�uBWp��\�;3_cw�J��$u^9sQ6���{z�&����#���㛟@��H������V5[I�]�р��<���v7ʤx
�k�4 �IQ̕��s�TP����̑�)��)��������K��_�yV��Zߐ�TlI�lJ����|��ә���P"�M|MD�VV��W�ůY�/��:<�E��y=q\�x:��];�Ț�u�W*}n>Dy5>�~��]%.�s�Ì�@�qI�t���v5R
�V�'P����qTE^x�yv��{����ޭ�����d���}���Ч�m� �N8�' ;���d�Թ����x�0�+����#�Ij�T!ל��0^Yx�,�B��L�kQ��\�KZPH��ߧ�v����y�����d_��h(+��u�fuS�Tˢ�dQi�Za�A�@TT�n�Q`!���&B?ՎA��既J͠�с�g>�ǁJQ��z ����͋!�5v��e�ʋ�?@us�η#��.=�d��"��e�f�v�*�:7R�tߞu�sS2p���W�oG�oR/�V#D����o�f��ۿm����u�Ymٖ]wY���x �G�_�>���IBN�7������Q� ��y%�X��ҁt���^t��|V�6P���ũi�2ns3����c�����6*���ſ@�i�JsX��2�Z����3��s/�Z�qn+��9��8�~�7�)_XY�Wn�eR�5�_c+$5h��(<�����
�eA%�?��P��[��P���D��ۅ������ ���6��*�܇����Gy���//Z݁��7�Q�^z!t���m�dQ�/�|hb"�b����0�T������/�p���]��JO�����JĆ�WR$�4��a�������뛈�)�!E*�^������"����*���a/|YY"^�"�7I�� ,5�ѬH�G�i��Kd����|��.���� Q�\K{A>�gq��h�i�!��������`���Z���g��G�?{��G�&ߥ�#�v��]���Wd��^��s[�OФΫN��S߈m}��G}ϸ_v���.��F�޾7@�~C�C0�f8S��v���I-[�lJ��&=�|���� ���4Qmݢ�!�A} cX�5�N�j�\N���8��"R7~hM*8漎��MY%��AJu�b��'��/Hd�?K��^���bQ�Q�;�IeN`�mt�(6 f��!4�༗���
�n����m���o�`s���_t|S��E[�Y�I/�[�#�k�Ӻ�X��*�&u�U쮋���w癧;�r%t����qWݔ��2��M�Pu6Hk���l�'X�Ps-�WYD�ܽ�v��ت{��%�yy��퐛�#��E8����Di%�tl�As�R"�Y[�̒X�	/�U7�wlHH�|��Q�"����)DMj#��߱�K�$/�(���z~�\& ���d�&�P�&/�@?u/��x�ԮP�Vs��U��� J
Y�Q����+uI �K"�bj���[E�kS3��ܶu��b*�U-B�Ϟ���-��H����aF�I�G\d�ډ�ɕ$���4�P��scAJ�Ǘ�hhg���;��=����W���oW���Sd��ݒ�;�Z�h
��W�Q'����k��� %�V7%�2]iJѺ�Z��� _-���.�ƞ|'�~2?��x��u��l�������~�N-���)aQ"�
�� ������(�=u)�z��ǟ	�#�C�v��͆d	�2eN�-�`P�-
$�œ"eM���W��V��/�=�u��5EW֡�X�[�
N�ߛ�Y����yߘj�`U�L>H�)�� ����Q}��*�|h����i)F����bGV���C�r�]l�:o�8�΅F>Ԑ����$���R��n�3ק����˶P_���]���[ep�c����e_�p��M���|�3��~��v�����di������s��D�ZnP��F]�0�pp&����*��_nw�٭��0\�'�Ȭ;*�+�p�n�<��U�j��zdl�VAz�C�����_��L��ѺeL_q��hî�sgi��mۡ�w�x	>O����2�!��c�] ��nt:u�섆$��,F�7��Z�LF�A�P��Sa>��Q]*�2g�vj��"�sm*�Bzz��i�W���ɫ�#���|��1��d���~���C��=���iw"W\�?�@9ͳ�����ښϽ�ZlXq�p���-B'��;����f?�ԣ��Oj����ͧ�M�U�q�U�C�;��R,I
`
�������/� Pv�wR���ԑ<;;�z�������!�5�����'$���;yB��w�s@�o~qY�h<�1��C#cn�[���e���!�G��P��f/]�3������B��9�{H�ޓ�W��d4�!��^u�#�JP��+������6`�w�՞q��e�ز�O�<�o�5�
��ᡐ��Q�	h۵k�"�O�|D;�ү^T�I��>v����aȾ�8s]pS+μ��m�}qВ�,iS�JǂJ�ƾݔ����SQf��QWI�M��}��D+�0�`�Cs#��%�)��d���e��m?�����#?jW.����l��yJ�RC�(y:�n �Tl-9R��@��-ԕf%�&�ר;�ȱ6����~�o|ݾ{�e���FB(���IzOX�[��T��Aj�.�C��7lW�K��)���@�!zX�9AH5�_卅�C
C�Ou5�&���~sh�f�$3_kv������+Ų���P���}9�-����D�2�?����	��
E��+�624�gb�[R��X��N#{u���x8��P�ݳ������?�i{�ٯ;hYPژ7�P|�T ������WT-M�%U��/.E<KARh�7	:�I3�o��V-��BE�������EV;�=��"�A�������st ��\���hY8D�8/uq��A<F��z�
���*ji���f3�3f��$�"w]���;t�|&c��4�Y\3�u����)��y��k`�'R��%�
'd�s�+&��Pg�&@A2�Gu�=����/u󳼰XGD��X��G�������xP���Yq/,u5K�96�%0��I�l�=U�C��:�sH1�BI$�kl>&|/���GѼvLg-��;O���D�i̹�޻�K�zޖ�!�ÆO}p���q�L�;���$�Q}��-D�d�y��'���3������[������A½�d��)N�2'tn
��S�L������МF�)yV������p0\"z�k��x�]��Ǐ��fFj��m����m�Ԧ5����;���;u��{i�#��N�{��Y��̬I����"��o~%5e5���	����Q�����jI�2.;o�a�.���О?���9z�N�:��%��29EB�;$�KFۍPCI����.�9�Ϛtz���c�� ��V]�X�a߀�}�g~-D.{)m���WJɩ�Ȋ���6ݑ]�ě��� ^�Q(v�E��ra�<z��ٳKO	�\p�rҁ·�bT"j�Z,'e�.��A��i��g�r��p���5�M�rumzN �X�js���=L�y�
��~/���J��xth8�^�Qp��/���[>�'"�;Վ�
�j�	`��z�ak|YD�ҵ��m$2E����!R��7��b�2�&4��S���9���
d�6�a���:h2lD��ɢzLс2N7B�����y-��
D�E�'u�>�� ��D��k�୭��W�L�>��m��*�̾H�j�X�SF��m"k(���д��zD4<��a��5�.��kJ��V"�{��2.��v��Q�C <���H�,�ԫ1�hc�z��}�� cΫ�#n���ޥ2�N�{��<u�����������bG��J�f
Pqp/Y�o$��L.]U�B�u.�Kbȗr�)]�.tڢ����.�۷���x�֩Mͻ�.�-���@Y��o�R���T�ܹ��@�>�
��E��+;�ݘ�(�-����s�	����ɕ7�U�5J� �T]��tW�)Jg%�t���h�S����κr#�c|̶����֚/AB�� �1�[��2Ks��>�H�k�Ў~U�˺��6���*-�L��R`�&Y��=��HP{r�m����&ʯ���o��BZ�tf�{ :��^:�f5DBߤ���E�ý�4��hR��L$�'=F�zA^��W5:f˽��F�d��!)�v��!��k���� �)�������|=�H~�~�Kdo�޽��*�QM #@&��S��
�9��V�����/-�������Dƒ��9�t-cM�Bn��ƅc���.2� 36��wt��'���؊��D�,�U5����Ч��Ї���v7Zg��d�ڏ,�-#`l�%΂td,�g���c��-D�ݚ�b�c�P������76="! ��M]��ou
��+K`�9�YZlX��_���q��X���z(�vCU���?˶�?[�>x��nIo��ӝ�V��u~]��N���~�R̬젤��r^��"wh.Jo�KL\��~&��e��r��˫��vc��g�of'�\��pWlَ�>n~}~jhG����U��K_�j�!9�g��f�f4���r[��T5�o��|��j�5ml(�T�ru|N�u�En�<[XY��� |�h�>���֨��)�����\��C���f+G�l��e9V�%r@�j�t��W��M@,�����>�P[)�lmiV#��f1h*w��S����4�s{en��ɪ�l��oJI�({J	���g5?�J"n/88X��-V���Ԭ�x�p c"DIZ�w�PZ����c�.�E��tS��y���R*.<��υ��Ru�w��ځ�QkM�z����Z�ЁN��G��� (��t�h"`�	`��9���>$;�o�Ϳ����"��v^�7�7|����'dK�}��b�0/;G�L
M
*�U_v��?�F�s��l�oמB1�̵)e]�������V+��:o>����ޅ��裏*#�wߌ�a����׀<(6��8�`�(��rA���������{u�|!�2�=sY������k�k'r��*�$��O��y���u?��3jʼx��?���0G��P `�L\�I��؟���1�_}��=
��kW�T0_Q�)�Z�Jh M$���O������#�((ύ{ ���+{��)ltT+*�R7��أ������ځ{�U���%��ך�q+eL��I���;��&�᎞9X����zKQ?J�$�U6{���<���ޚ��H�c7��\���c
��G�	���vB�Q�Ty�R��[Y��@��[�8򑵼mC�6�vţ-}��6��2m��XWB�a9W�S��l�v����T�"��m�X��y���U�|yB�CpFɋ"��{l����(FJ��?��3x�`�Ff¾ِ &0�kl�Vѡ����/DʚZ࿣�q9�Rg�u�CQ��9�k5
ƫ��n�jU���z]����L���/Md��D����!�SVb�~'jA�5lx�����Q���i6CS��ny]��8)�ҽ�\R/�D &�qtl\�nD(�[r �?4��_𚊖�9XԀg�|B}H ��1�GI"���a�Xx\iu����rDu�S���
:��WȽax��I�G��
i����ۈu(���"-.�E^����>��}���7>�&;��a[y�娓�ۘ��M����4]��C��H>/bSJ�FJt�&�0�m�Z{��|�Q��� `՞�2Zx}�Uů{mq^e-~M��h<ZH�QSR��:��NI�3�5���.OOؾ��(�䆫��h`D�����ʶ�0+�u�N[�[RAu�X$e0#(�G�q�F��)kp")�p�I�Ђ_C�޴�}ؾ�ܷl��i�g`�Vf/�����>m�s�v��)��q%s��ǁ�ֽo葐�at�kk~�V���	�ڬ�C�(B�!N��;�e���g}��~�9�^���������}�ݩ���J��}����c�w��b��u�U�F�����x��o�����NOm�P$��KtW���!��}����-��I��m�	�D�]��b�$�dK�� ���F]YuR�j�?s��쨝�Zj9i.�y�p-�����q(���"8t���v�ʤݱs���v`�[��Q��S���yEH�0acuh8�ؽ�rM)W6�B�]��$g�nk�m��=��ӓ���+�)
[����=�7�lS��o
��{����������_�'Nv���J�;;"�S�� �iW���U��x���p]�pV�ؾ��2l�w߭{XV�����d�@r���{�[<��>2/8.��yg�i��=P��4�s�[��ɴr���D�}��R�D8q�a�����^���)*�[���dkٛ�\�oHu����:�������퀑k&bHT�́8N���� ���F�&d�V}O�Q0���ed|Lcɽr��C<�%�?S��lc��5<g"��[9�����]?v{ii)֬SS^��u|��?�qTF��3�/���kU�$����P(�D���ҥ2.��i������n�;uw���sj9��B|�o�4Å��}m����Uʺ���^��f1��yM+�I �m��,��ģ��wnT3>Ȏ���� *�O�^-?&哮��Խ()* b'4�t/�Bj�(�J�4J���dw�u��ZV�uO��P�����*�)��?�����r!�f�/���![Z�w#J�<'�M�z�(��x��^.1���@S>4��#�ƈb�+`�KF�ڤ{N���O�c����S���s�ܙ�Vl����Zp���u*H_��Đ���5:����	X�&z���i�j�˧i�St1��åG;D��7_l�_S3Ih�	n"�m�|���J�0Ģ�E6�����w�n��U5��ɷB;"�p�I&j|��E
< j"�PZ��r�)i|��"J8��5�fhpX�Hj_�?P����e����/���4�"�s"si	"���H��5q6�w #�)V�r��E��a7� U��p�Й����f�0���������{I0��},e��z�!4���/�I%��u��ͤ6����9:����h]P㬀��B�YE����qM@fbzƞ��v���Rq�;()�۪=ju���Y��n�����ꜵ��DkB�a'6�!s�F��������˟�u����;�f=fJ>�|�_������G�����oz�~��?c_����� ���cm#�h�ک�E���G>�"Yj�}~,�܀��w����e���?�ðh[+M{��m�o���9X�9X��6a��s��j�F��_U)/�Y�Cv 5s��E��n�a_O��(�Dg���%�.ϴ�
�0cgO^��݃���|�}���g-[o�������k��^:z���?�W6�N�����	�ើ^���f�_2�>(iE�C���t~>�TE�s& �\]�7�����ǭ�k ���������!~�r�Y�P�:9��>�aݦ|��[zG�$�X�Y����M�����1�+�m�nL>�s>���ۏ�뭶e����><���>J�ZA���_��,�
P��3:a	$��9 wn|PN��;�Y�V�����ew,��u|]���7<j[�v�c��-���J
��ԠR&I�к�p��ksg�:�1`"��BN��uW���uq睷ٯ}����o|C�ru}�܊��@$��H����c�|LM^S�h�m��ȄJ� �޽�Q��-˂]�F�t�dC�2�������e?!�ý�r޻o��(� �P��V��,ʾ4�㵊�-,��s��_r߻��*�T�>Ҕ-�AEY:�Ѭ*�E�)� I�;�pWu�C��LP�r%�V���?a�K~]W4���v��U�"��'K��q�.�q"�D�����FFU�t]Tp}���X����`�˕�Ad��l�6.FƅƝ�a�|�>b�|�;CW�Ԥ�@���z*���#ZG��(RB@�wK�
!@�>%���+�m�zH /S����S)������v��i�m�k���3ЯR�Tj�p�U]˚ӝ�%�\�4w�#��1/D~glƷ�m�z��SL~ �l���/�dV�43�S^	�u��K2�:�6��6�0"�r�*�u'.OڋGN�۞|��aQP�`G��y�^�/pő�k��&<oHI��,f�7@+�L�)�g���o ~RnAKf�ݍ�v����u,I1	&R�D� 7x7P� v����?�w�{N �A'J�D
��3����S��DϢ��έ��ױ���/@�@i6�����[UGB��n�J��eH����`2���w��WcN�/�Z��U!JE����5� )���2��%<'�v,��l�Ww��%[tc���C�Q.���:���W+=]�$��j�����cGC��~/�3�/��x{IcT���7���3$�o
H�l�7����z7b�B-N�?���^��S�J�_��w��(�X ������{��z�R��Z�azl�I��.��Q���_�5��k�A�ڝV�Mc���L��^E�r]=ܰ��Y�@[oa��oX�=�����g����T���WWT|�⇭�r_��nw��gSn�:�]-:s�Z��ku�Ulya͞��^{�[���-cv��p� P.*}H�y���>�۽���سݞ~�.&Վ�����t��S]��v+�ۊ��t���<v��۽�O�}����ڻ~����%L��o�!��\����ū6��lnj�� �ۅ��ɎU��� j���>��o��Hg����t�T��m��{�}�a{˟{��.�����.]Xh���>w��|��:�2�Ͷ�n���K�A�ȑmY`1H��V���spe�4�d�����;�!�� �{���كwmsgҁ�ۨqꜗ�c>߫Ҍ�c[(��׬����E�����`a�;{��Q;}��8ëHD��"j7>��m���-ۜQR�
����\�c�Ϲ���gK(��Y\w�5��ڠϓޮ�n�U����������|�Z�̮^�(ʣ��Nټ�ȳ�'ltx�.��];z�n۷K�>}t�Gz��2��f qV�H��3\�i_�Ε��N��9����  ��IDAT;i?���'?i�����4kK�M��e�zuý`G � �Rߒ^KI�SǂzJ(Z�];w�Z����%>X�3�x�q�^�/���oJ��<jG�K�B|h��U�g}A�s�}��0|�SM7{�]�nO�=�ٻ����S;wmU�3���=�m9�\#����p�Le, Mu,��gҔH���W�棣K���O����^R�\����_������!��}�鐵�K��������s�R3��y>Ԥ��8������G�/�����������*֩F� �jyDQ��}��+v���u�����;z���/�w�/|����Ts \'�?5���v'�{���_I�E��&[�]���\SL�b-i3:ɛ���J}8˂�l�/���Z5�S����7��$����NM�p���v#�u6�T�L�'Bֽ��K/����ط[��p6l:�-�w���^�6z]��>q	��=��!�\�ٌ5��A����_"�-�Nlt�_���wqhoo�z:<o�����?&-������}�_-����bj3����(������zh�MB8z��ih&#�;�"�㽄�yN ����>{JD�ը�9���_hXa2R��u|�]L�=�9���xѭLSQ;舒�P�fzR ��gC��_����sm�:���slC
'�l�{����ˬ)<��|��:��'o�ԘR�׆QmEY?4�S=cA\�-u�j�ga�tPK8��18��c�����Oػ~�]��c��ۙ�eP����՚gI�3 Ŭ�Cs�MS���1Q<F��qn��yo�R1�\�SS�6vw�f�r���)�����}I����(�� $�S�<�pD��̑�RSÊc���"�a]'��@��Ⱦ۬��qg�v�Z��2�K˽�\U��c�!�6ܙ�k�"�a�� _#P\n$��'��n�̢g��r��:����)��/�;�.�l�������:�{W{�k�=e��3h��畮lv����%��m�lt��y��
�)��z2+hl�ei��E�� �D$�C�^{�G��/#
x��;v⤝�z�
��&��;�u�<t�N��t;��y>���Ȯ�1�r!�߃W_�G;T��rd��k��2�GYg8D׮��E��V��k4m��`���]w���862dC�)(�sQX��-[�mt��._��<Z&��$� 
�My��S� �c,�fuGϯ��-���_�[�m��[�TU.�O�����,��>�JY��+`�TX���S�q(�T!�ld�<�^�"f�]���)��\Xo�=s����ݲS�A^����;�Q�Q)Ih�
�|��**H�_�H`Q��ѱݡ؟����ߔz�W����ȸ+��v�ש1�7z)ά=�+�CL(�	u�kk��j�;wV����{�9 Mg �7=�F;t落r���_s�K�k�~]uܨgQbt�mM��A�CDr�A�n�����9.F��_ ��ٳz�b�q]{��⬈�x�.n��E���J@���Z���2�k�`$�z����kJ��[�q[]V-7ӌ)a�N"¡���k8D�,*�%
"�Jf3�>���X5�u. �J�q/����5 ;�워��o���w���c��y$��4'n�u8L�V7e>�"�N�$�ɬX����u�l�Xcm٧h��{Վ_�f�Ճ6��I��_u3�:�N7@�9��ۚ��k����WK8����wT$�Y���BMP�:��E��z���)]�Kб�'T��k�]���&b���lB���j���`x���?������Ě�N���n���6$r�g��T�IC̾=���>��3�_5 �T�F�H$��;�U/`��q3Af���8��4-��М����h(����quF��o�*��)��f�Z����R*+tږ|2���j,������Fqs�"`����jd|��;�^5��(ޓ��Yd*"�Lh:�6�=�����5'���B��n��=،�΂"o��ރ��b�̒FA�,��p��,��n3��g��6pJ���`dI)�e��#�_\�;~���/�<R�pa�C�G���I��b�8����!�\Z�.f�W� �!I-$)ku�j�5����E��4R:!P���ki��ş���:�%]ro>�F&��D����z(���.-���Z�r��{M�9(_N:H��?��!T8�k�--���H���uS�h�"�� oJ$E\]&��j�T�s�^�OV�%H�t��;�srx7Z�h]�\�#���_^g۠mh��������?���L�SjG�������`_��foz��HAi�IB3s��;0jM��_�������!��Ӷuɻ��YG�1�4{ �� �Z�q'*?�v�L
���-���:M�]�;v��8jCż�:|�>�۟��}�K�$��s-+T$�Xtп�Bidؿ���Gr`4�UD�V�0�bG�]؅n�ߓ�����pi�>����ݶk\|�5��O>�ݻ�6��]������W��˶��hO��	�>2hg_9jo}�����u4$MJd/W��zF�R ��us����\�M��h�d^�N��;��x����[~����>Ss�HS��,�E�ulBVok�V�4F��4U��b1��&jUD�p����mlKAL	�D�s�̞�@����[��Z1��E� ۊ,-���-3*�M=���k�I/�)tl����=����H]��}�/�3�ц�T�7��ơFW�}{����	��� �F�.�Y����> {�@�Ͷ�,_�C+��A�ON���괫ڷ��t0N�"�~M Z@SPe١�2�\D� M{v�R��,|�n_(Iz𡇴?PY�����x�ĉ@�-Əye�HuS���M�)�,ƌNn��7X� �Yt���4����O��s.D� Z�[U�>u�������pW�ki)У1��������^e�`� �n�M�YL#�ޑ�z���;�Q����{Y�쾦���R��kV�uIT���������Z���[��@�;�t*�������Ő0@P+I8�}:�u��47�e�<��>!/W.��{��HS@�Q ����nm��r��m��:�N4*�S1��s��G�I�r�(WW�v�ʄ=��/�J�Z�g�iJ��\��3�]nK7U�u�V6��nYC�$����I��:��z4Yj�Ѱި�J�R�N��;h���ZY�YL��b���d�����#=l��jϻG��3��x+,��>�����F¤�Z$.?��Ξ;�t@�{Ȑ��5A�}�A!jsBڊ�JJ��$�d�� �Z��HU_��'��B�k��/YS]!��d���F3E3���.�A�A?8P��\��:"Ɓ�]̡nOrN���#*P_\Ҡ!`�>a�(�z7�0�G~,6ujV0J99�
�}�u�U���Jc���ZP�`�M��.7��߱)a��s���K!��ы���=�~�;��(��f����D�{i�F4^�@�$<�T�Ab�MOMj��=_uZ��t
sB48|V3�}OOQ)��o}���lJ���r�� j�_9.���Ј���>���]%����-RT BaO�-�z�D�`2!��w相��= �5?�d�e��h��Sq�B��*�V��*3��He��[�yg�7Ϯ�j�숚�hZ�v�g'M%��{ƍ���ؔoJ�>&[�ﲡ�m�Y"�o&=�]�4�\'d-��(^�~��MB
�D[�NMҝ�3M�6��w�q���SRvg՝��c�햝R�N����_�/�Vv0�V*�z�f[����nC|���=j+���'#�Xɭ=D4z�P9"��kt�bmU�H����5;;=o|���\�6i���cO>���ˎ}�?g��f_����C�-ߨ����8����7+꼎��������l�9r��@��ې�˅Z����e��;��g������sV����~�Rq;����U�-��Nϥ�9�����)����z夗KU-��7�v~ƪ�q�8Z��,���M.]�XW{l%^��(3(��`�7ST�[_�@��h����M��r�"�{qN�?�3?mO�i��,�5K� iZl.v�9�c+
<�Ā��r�ۜ�زՁ�Ve� ��G����*�u5.������|u�N�:-;��AZ�ssv��a;qꌾ�g�٩�R��^��1��^��f2uʣ���Љɫ���E�C��n��6q@RF�iYm;z��_˄��5�p���צô�gp}~Q�yRDTJT.
�s-�ɚ�lB4;	h�v���f���X�ؑe�9�6Q���%߃�|��~5�^8^ײu�X�ݭ�����?�w��~��
dL^��B�l�xH�bh��`�f�� p����7�ۮ~�V�\����f��Dj��9�q;y��U�ғ�u�Q�DN�xZ�Y ��h�ls�H��.�D��"�F��C#��0��g���fCͦrgSk��C��nQ80��vn�vCmR7�xS>tOߐͺ;x��E��_�>7N%�u-�#��z�
�N'���h���h
i��W�i�%��s)5�{6�*@�)Ⱥ�oY�c�}�h|� 
�lH�ƽ#"}��.����_��_���[�e���gD	�<�����g�|O �H$�5�������z�,<'&>���Z�K깨&�u}�1�?;x��al��(e�nS^����`<�I�e�;�ݶ́ݔΙ<8��Dh.j��$x�%�E�d*0�<as�( h��=$i�P�T覡Y�t��g2R
5�����o%��߸�ϝ��ג
ZRSP�����w��ȵ$���V�����������;0R'��}��+��K����h�4GBD0#zZ�?�1RT�M�;H�E �rm|Ѹ��Iʥ�-1
��ư�C1;S��Om`о��o���X�o��T�V�ޛK��~MŜ�[�z�r!�,MQ��C��D�j����>m�k;�z�X�����s�{���;�Y-�D�l8�,��z)c4��Z����"T1
���&u��sŪ-�i,)��.��Yۿ$mC�
�.��ƪ��"��u�B�(�?�lٸ���������)t���c˜�um����2?7+g��ԫ{]���ȭ!�������׌om�m�s���|;>�)��Q"i�4R�V﬉�Ϟs(z��lA��X�\�=��8\v����I����疏[���ײ?�m۵o�U�
��ۖ�!�V��󗃬!��Mݑ�:��=7>Mm��T��R�E��^9ew�ն�2��L�;�is�b{��"��<&����t24��r'&�2�����с&��ڶٹ�v��u�t�5石���hw���:���UJ'�3Ss��H�f����� R=�8�b'.ٌw���`A4M�k%�^����!ʕ��i"��KҴ�Q ?�޽G�H4Y�������k68�/�F�I�F#{26�E3 ��������싙$ҵТ�:p����~�WDC��@����b�@�H��Ŷ��LT;�29uI5�M5�u�]0&�H� KI,!5��R��]]��E��"�g2Ma�,&�1�=�8u�=g(�G2s��Q�Bmu���F�+W/u){�1��#��C
$������H�o`���C�)���u�U	��yn�{��N�\m�Ԥ-��̝��3���_��5�n�2�E$_��/ �j֙�;��r����\\�I�2�d<�!v��. I��ӪE����Q�"��Ь[���H��f )���~{��i�66l;��j�ҍ(��FI=bD�x�����\�cڌ�t���Ҕ��j^x8t5���B�~�jm�ߨ�2�qw�;T
��?�P�G��	�B[X�}���O����?�'h_���
��o7��8Y�;�L�%u��K�D,ޤ;) k0��|�JQĘ��w %B����Jw��%	�V�T�RT�5Ţ�0Mf�����w�!�c;���깳�����9�/�q}�@y!�k1h���7����I���+0����>���m���&�����DF��� �$�^�A,���t3*>� ��}`v�x������WcC:f���V��)b�	��"�nY..�D�މu&aN�K��$�j���A�)5L�  ��Pn��p�
��X�c@PQ�
���]���o�tĦ�-���Q���hK�IS�a��wu����ْZ���cA)o+YӖ[+۳g�}��9:�l����}�.�ܨ�L�9)��=�B"���$��9�9d�@������uR�5Ք��qoB�@M_��4�yޝv#D�,��Ey����e�ƮI���H])
��y�7�����}"�M9	�*�DW�[�Th��Q��ʀ�i���*au��^�����"Y
0b�x�#���`f=�����D����R���EY/���;ܧ��K�uKe�F_Ͼy3>0M��5��R'Bf����=k����8��u@I�;u}�pޔzk{�AO����~ �s��uj&lf~�^t�v�'���yȣ։��zI��oR�ؼ���5�D���7�}����Ҋ 6ه�ЀY��>�{�ח�������l���"�Y��y��z�i�
�c�}}�(��ҩ��ܼ5t�����Y�nñE ���:��?��?ssV�ée :�����k�lIpx�X�`K�"îOLM؄;�;���s;�&%�	�����0��]�w�;2;�G���fl3�LMc���#j]����ԭ۷���J9�ļ��.]�z#�9���a�Ϝ��&��8J�LJ���-��<==�=7d��0 �r�sjMr�����w��$��Z�����3�c$8�}2��@p����#�_�]��aums=�"p.�Ӱ'��R�A�$��X�={J�+�@�{"��wkn�� ���]s'x5�ؗ��9�|d�J,շ����@/᪛zq_U���Q��)fzs��y3단�65�}p��d��
�x�����,��n���x��Ǭ��CSgdmh�^<z�v��c���,��CǖM�\h�>����U�j���8��Vm��4�U��w�� H�=�B�J֏�wJ='P�"��;t�]� bX�xU�f����o|�v��
p��cnf�ہ[�rC��F�pj�~5�Dfy@���':�Ddn-zOI� ��Ib�VS�/G!����l�E���)*����I{� ;��L�d��_���B,$ �$H�"ŝ�i��B�Z,[c�����{�v�DLL�����c;f��v�L��n��˶H��BJ�Dqw$ b��W��e��;��{� R�'�BU��/����;߇�$"U���4>�f��@GO]Ĩxp>������;q�	{�9�=��z�$�1�A6x�!�9d�s��Bƪ#���e˶RnI�T Mb�@[ ���3�x=���^w9��QY7p�M���cN�	j�z�A����M���;x]Ǐ~�NH�_�.0�2M�^#�A貊^�����`ǩ� �Ÿ�9��E0�,"W���6k̆�[�Ma��0�d|Q.�W4�Ͱ(Ͻ�=wY��(˅-j�$놃M`�<"���U�HÌ�
�y�n���Q��M�8!��{�n)��yݼ/���Vvm6Vd�������1���ԑ�GU�ݕ�%��y�� �Zs�Ў�7���5��P�~�� ���A��} ��~)Y��cC�NJ�Բ�ǖQ�H\��kZ��}�����Χ:n�V�X?�'�h�E�y����q�:t�����:&K2�q�T6hp�`<):�#a��gCD�zlh��q��eXL�G�)*��64ƬHMmV��]6?�٩49J�M����SWJ:G\8wF��n!W�+E����K�qӟ-[�at>���A�cY>���?��!�:V�ﺍR�eu�M:��6�F]븓���v]�T0�<��~kd���dE��Ƌ��y;4���e�*��xl�L'��ɠ��b�����+.�������{F0�sjP��c��p�ppΫ�����կʽ��'���c�o}����cc㴝�U[q������fcP��MB*MKLL�˘��M�gda�2�)oUy�`���֣�XU�j.c:.P��9X�W[e��'�h��G�_����s�rT�|XE �4~՛��fqai�v�6�?!�Z�-�$��+�]��ubײ�8�[u."����u_�f�ef����I�8�K�}�l����\���Ǚل��;���t�AW�5/<��������t�MtN������e�)����D� �^������#�'5��܏M�Q��NC��D֠<|[�|�$'/,���+婍��d�Z�}��?��$�o_3���Y�r�����S�Z�R��t��5
��≘�4[�������%�p����|�����2�!%�N^8'O��%ׇ��6�C���K���FY�h���ȁ���1Z��R]�e�3�@� �EcvG�WD�>O�Ę���O�c1x��q����fL\�N��#���֐��|�1\\������N��^����{y����Q�H/�]\wQ_^����z��#X�p,0�]Q��K���Ҋ�Y��1Ny�K؈���`SB� %��'�s�Qޮ��+�Ӻ��]^d��h4�j��i|���
]�C�zaȖu�CQ��~�1�7��Ɣd���a<���؂� ���_(�W+&i85���;��!��#G1�?ݜ�G�x^tf�:~R.���Y���I����	�~q����/ɭ����y�y>{�7�p#QH]a��:-�{%퍧�H���;�~S!�51�l�itt"��r�$�`71"V�\*!����#�	|f�g�R'A�3K�:�
U�sey��w�w�J�����nk�H�i�d� �^�eagZPp&�>��2*�@���r��E�f��{���{���u�R8��U����+�y�:���t�[k���J.��{��+5Qu�<K�8gk��,�:�L-#R�]��۔���Ay��b\��F���+$�}�W���T����R�0���w���
����k�i����Iu���s*Ɂ�{��ݻ$�u�,�����N��B]I:0�ƊW�2Br�#j�4V�9l��7%1^T<��M� �����J��G�q�c\7��+zuRP�m����鹷��A�ywq^J�T:צ��}�[e���v��ws��VuS���r�l����ێ���L�����p~{U,v41 �Z,P���w��kw��ȰTFЭ�!ޜ���J��sTQ������	�h��NMLȤ2�u��]��ĕ�tci��#����w?����M��� ��AD�)u���.o\G'6,r��p�(��G��������)p�HJ�a�x�)l�(���`����Q����B8,gN���8�8�*8��!�qaVË�1�ټ�N5���Mip'����F�
���h[������M�0aR{p��<��������� ��R���1f�@f�,"Fd*�C#���W��ʥK��`��;����c� �^&B�qE�<؇"6���ևAO?�k#Y��{:��ã_�g��p��c�N��Y_��YQk��}ƾ���[��}�r�k�ɝd��2�"�F�𰰝�Fw���j.*YE��C��l�:�ż����n�9�`�
e�[jw
�,�Ry���e����a?�d%v�&"R_]���c}�UVB�^%{!g�9�	.�%9����FZ[^�ΕS��A�N7�#;�l�$��dy�.���}uע�>bb��9(��[�wu�L�S��ZRgg�J&�f��҈sV�3��tм�$�R�(��T��Dy��bja����~��z��On�������&��,(�x�n��x�7醊�շ5�����ϙ9��6�a�##��ƣMz�k�|��\�}ibм4��IQJI*B8� p#�A�`j83�slq�MP� ��CD�#�;,�C�=�sC6(�����A��%}�dM7�<�P��c�63�x-�Q�i>g� d����>���ͬρ?�"��W�`�!�������G�z@��%ٿ���׾&w�qG����h�88��bDxb}���-aVf&n5�e?@F�	�Xe�*2I?\��$8r ��c]��Ց5�"�-��c�WmP�5�W�"W�ʙ��γ?����X$�<CX��%?�K��C�*�5t`�C:�g�9��/�i�פ��럾�=��O�77�_��gd���wrr�t����\쨁?r��u�nF��*$戥.3K̩/;3���y�bd`�1dn�s�,5������V�j��6G����ʧ>�SAVg/Ȣ5<_G�õ�\E��W$�E��8;S�W��P)�n��;v�W~�����dD/qK�A�3�E>��_�:71'&�GL"�A r������?��xNF7]#%u6��T�@�(ԱR���D�7zr\ޙ���X�OX��!�7�r�|]��?yEFF7�ѿe�.9p�u�V�kT��<�=�k�,����ܹ�z��
š��+Xd�u���YM+j�_U���â�o%�S�"��q͒6Oc�3�p���@U�7g6���Y����L�r��~�yY���i��ZC��T'5�c��㮋�����u�vӮxf�(�+6 `̢ �T{�e�X4��2�)]�;�S���H{�;��<�FGt����}�v�78?������f���]G��˯�=�$ ��`/A6���o0�r�G�#��,P��\�p�I�0�(7#����@j}��4���$$��%��3�Dz��w!��0�Gd7�CV!^U���	�x�t���R����=���2m'�{a��H����s<p����^�\&U��
�Q��2���Lɢ`U��4�<�O?�ρ,!�J��S5��y����H]����b��p ���-�=����!�C3�L�+R�>�<�����Q�sz�V�y��8;�}XC�胎��<�$�Uvrnަ���,M�,n�����1���U��FF�s|�a�n@L]�;;�|wNf]6��{�8=�'1R�d7F9'�0�g�l�(kKyy��)r:�~�6ׅS[�LrϢ+C@��]>��t��2p; �y��ur��E�I�A���$������������.]Hp�`�:��:G�-xNL���~�xA�� ��;��^y���o���IލHN.'���� ���C�0�8�0,����E9r�p��9p����8���g�/�##֐����0R�6�-���J�>6�!pZh�@	�_F7�\��bp�|���aM�.�����/�3�2J1`����T���:�lNV��¸��%���((��1�5�{a@6m����ss��PZF@a��Pr�[�W[qϏ]����"�0�A?���<(��ę��<g��`a�æTw�#fe�y�F�YDmg:2Q_k�u�����2���{��X.՚�ҍ����p}正�j��hZ%��wp�������KQ�к�jK���䞏��l�t�*}��
^Z����έړ��7�#�~�9i��:(�R`�d����a7镞]�B��$X.��oqU6�e��>#�6�ImiV7�	:�ؤ斖�֨˝�ܭ����wE��vV�����T6�݊>�5[�r}Xw�����~��ɻ���y�ΞPGc�O��P,;o�-����DJ��XW�ǁ��ʣ�|T�~�M�GeT��Ĭa'��]�q_O2�ڣGJ�K�$�u,m��4!����Қ�}�l�f�T����%7��'��1��Fԡj��$ұ{���=/�D
#CT6�3��Z�T`��Os9�2�۾�j{��B6L�ڱ���q�ܰC6�U�	�`�{d�N�c|�JSU�� m0#[�?r�`����s���o�	
�U�6��:�o:��W�u�u��gc:H2��g	��)�A��C�JҰo��9s�}�!���7�tݾ��/��Ȋ�*t�^�7��o���ʓ?��<�
����쐩믧��ii`w�G��K�UM[,F2���%}�#$_^Ӡvv'W�8��VPn�8
6�<�7�P��-���ϗ�I����7���Z6��:����2c�|�����E n]�����{���Ö�I5ͨجr��ڜ5��[�A�D�8/Id����dJ�B`\�j۱`Bbibb�YP�#p��Y���g����u]�'|��7t�s�?̬�o��z���>A����G�<_�{�MKD4u�j]!.���5	��O�;%GN�1!�<�����s:�K�
IFQu���a֠�U����ɒ��+�=*,�w_3K�ԺE�L%��_T9Q%�j���s�
a_�Y� ~t� 0&��udb9���55$�l����qfPb�`�\���F<���)~��7)��iӱ5�B�2����K\�c,����$�0�S+��]=0�4���%(�:�N�?�]s:�8*�����C�I:��Pu���{����<�������S�����cH��:��5�P�å� �Rp��!�H���"��MB3��I�&t�'8�p����t��a��z?�530���xE���e��F�m��8��p���3;�L$��WA ���4q��%zo��:��07�B���CI�Mc�{��pyVN�<�2�?�_0�p=�%���8�wA�_��#��lY���oI�7����+�9���:?��<���Q Ŕ�k�	��J���.ZԹ04:&s����c�O�����g�ᒁ�ݵ|�
JF��*�A���^fJ��aS�!��X7��)y��{�W:O�K_�ͪ�j����dvnU�7TYn�������:���f�2�Nne��?1�����;�#؜��b��|��U~�s�@���j����ם�8Oz��礩NxI?6�[�z�EC�f�I�lp�kk2�]�FB|h��&F�ء�嶛�H��(��k�F'(xQ�5ȏ��a�S]A2��lzlB�8���=s�� �ڪ44 wm��8��g����\�w�?��5#�l,ݰ(�:�t-������#rݶ)I��2<�TG�,�Nm�(�wJ��O�9t��m�3�C���L@p�#���?V=��`��3ev�%���v�]23��MDij0�L2,��G���'�lSw�~\���|
4�PVGCݘ:̣ӛ([z���I+�[n����yF�{����
���hG�����K��V���f�gl�'J�[���Go�>��Cr��?�F|��k����O�8I{�k��N���K^(茡r��Nl2�����-�ѕ�>�,��S���l�Q�i|&J %'��Q���ĸ|���e$ٰu%6WZW7 �|�sS-E;�s�	2��:)?M�O�"H&lݲ�P-d���0Hl�⇽����,�����7���DFYH(������"���67�Hd�1��#����qM�>TR�Vn�DCoM�Z�p��s�ȶ�B2f��
 �x(Fu�85[]�h`�m�䙗ސ�U�e�*0�`؛vf��^��f�#�sR_s#�p$H��> N�Ă�&�Gn|bK���b�,9�"W��'.�F	ڻQ�N`��N�l�1��04(�%Ǝ��`�x��Ey��w�r��uzB����� t"��u�!��݌���f�+� ��l��p���K(-��?TI]�R�0�E�Ŋ�q��E��v�A���e�',�N�.��|�Y���yY�[i�֬1B�w����/<�	��o}K�x�	�r�V�8�V����j
rӾ����2��HrS,fDY�bY!��.cL�)jj4 0&���w�a�"�S�TV��$�_Z`�ѓ�sс��h�=m,Q :���r���X ����Ν�XR������X��C��ɒF�0 XX��5��:r�����$� �$��!z�h�rP֝�1��O�fW��:�_��^�������q\�slX�uءЕ���X7vgf[�(�c�H�S ���Ɍqah� ˨�P�\Tp<�(�S�9 �nS��yf�S5��T��/��t�ι���c�gI��C�:�8/�=��,+U�H�=�:(aW�r+��2�� ��o?N/u�~�U��%�	���\]�G�����pB����:�����r��9���
���iu�&v]+h�ʕ%5,��҂��zu��7(��Y	<�R��<Ʋ�'E����i�lz��b�P�X����JC��ac�'���2\&�x�jM���E�ǋ�8���������_�y���z'-��x���ݻv�]ԯ��T��5�ϴ�s�GA����E2�:KZ�.K%�Cn�]�/2�>� �ևaH��k��u�P���2����X��*����Z&��l�ˁ���5;vʙ���Yp�M��o��g%u��:\d7z�d0�Z֗���Qٌ"-Q/�*|NS�t���\	4�Xe��()LH�x���I[&�u~��"�J�k��.�z�f�͛6��wyq�{�q[�X�Dת��}U���ݴ��'c$���-+�U3���^��b?$l�ߠg�0
�ѸgV+�{wc�&N��L�o@Df��?K��^x�#xqa?�n�q��1�;'��oh���%b�!��=����6R�u���+�b?6��qBL{ٱJ����:]��E���hкŮ���KL��yo�����^������l$�2���.\d62����h@Zb�{�t�FC�{9yꤌ���������l�\���B��e��pU���<�����m[�7��u���?Mmk�G\�x^��F���3�@1La��ǬO��$�1�C�������l���1V^Y*v��^d�Q�*S1�!+��ԥ�����v��xT�;� !��ٶ��^$%p�޸{�p�2���;�+8��c���I-[9;�9k��^�(Ȩ�<$���\�D2I(�xe���Lؗ��a{��M�)�Ey��!���J���xR7�7��!����2^�pKrt/�n$���M\x���+�ĉ�7������D�s謄��
99[��B.�^D�u��='WϫzF䋃^x�8��J�x='�ð ̻{�n��?�yH��w�}WN�>%/��#A8c���]�x��� �6��F@�k�@�Y8,��i��:|��9���S��L��9��PrN�3�↓�#c~>��	]�2z����zI ��:�(���Z9w�,1��TW`	RvD�8��}S���xڛ�������zݲ� m][�3	���7�&�׮s���lAx�\�9�'�g �'�F�y���Rf���]�����3��EA�(�aQ��з��z&!'W��+�!��鰮EdꉕdI�����)9siN�B���n�6���0�:����:���v��)c��	���l8����Ko�!�9��~B�m^ʺ	�S2{�,�	�atWWwTʓb'F��wN�k�2k�릦q�o��%5�u�~��E	o�A▽��g�}^7�������Ę�LN�̖��DrqnA�l�P�Y�C:`\�c���=tܰ���g�a=y^�F�.���'��'�%74��L��y��]����*��8VG��-l^�&͕�L䷐�&�LO�K����t�3�l8��Z���f?�3�#����٣G���ʫ/?�r������Ј��1*�O��BN0��66�6 9�!F�c@��e=��"�R��.�Ӻa�~(��{?�^�d�XP�)�	��Tf8[M("f��s��EW/b>�gn~Y����Z�K�����ã'N�Y��n�ϵ�&`�@����#}M4x ;��`'�>ȗ�q��(�c?�
����l�~���GF�����O~R����F �$-ǌ,�&��F��zXfu,=^�n�����.l2���P&0�!{����,�5���8�/��(�#y�F�Eg�%f�	�i��h|aܰ?ў�^M�ku��Dd}71�hp}U׀9�=׏�ރςF5*h�����ľ�;w�W������I�BO�S����G�Jm]���߳����UBE��M�ֲ�pd��ۤ�L����*��j�V��������uK��"0���}.���`p������;p�mO��&<�bb�VE��'�ʺ�-���ޏ_��Fϩ�N�г��@$N��[�6d��G�%��w#�������6��A�Sdo�Mus4�~_�6��n�-c:��:腜~~�:=l t�F��sj|��ǔ�ۂ�3T��a"@u���#b���X�/4��&K�9W��Q�9�m
&/�zt|���k��i�۷�s�='G�׼��k�ڶc3t(C�@:���1�{MK�΃E�5'K��Ř�ME��.��'�."�T�:�}�%�Uq��/Q׺�l$���z�\ #�
,R,r ���z'ecS2AyD��q=(���:�H��0-	�g ����w�)�]�ۤ��jYSN�a��zbi&�S�s
���wӶ[�0l�Ӧ������#0���7�����rl��:�D���V �!#g6�EF�L�(2��Yb��5E4�������˺��\d�< .4�b��u��p4>c���=f�7$�H�(�c7�'���ٓ�V�\���pT�;t�;�@>��Z��λ��C�ʫ���轕���v��p�}M�7Kl#�;��F3�TiP'gny��=(��ߓ����=sQ��ay��qɍTd�����_��LV��SR�r�+㛆��la��Siq�.'90�:��*jp	Gq#x%wm�{�O�>zL�>yN"��:�jIXVB�gt� 7�Q�ˁ�r�%ӥ�v�,�F�q@y��m&׳]u���Հ=�'���X MY`˺T��ח�c��$�%<Ǯ4VV���+�@{hbJ���FG�L6д0b4�[>C�S�Y�s�|꿦��'� q�R!K�ds�̟n����.\�#'�ʾ��б/%�-�Σ��35��4[��28�Sf�Pq6�pZZ�Y�ذ�JU��BcUV���Ҿ�{e�4����ȸː��}+��id��{�
?��a��-��D�@U��{�"�ڛ��%�<��<�j��'R%nYv�vxaP-�V1�J[V�k���c���8p@��Dfp
0�� `xl�_���:c�L'F�'\�x<�8nR���h���L���� �_�9���jS�A��c�o���g�fP��bߠ�Z7�8�������F�1�$XX��`�J���؏Ο?���96n�����a�v��=뮞�R=�fk~���nf�b;xƘVG0�5�6� ��=��� �Oqr~��+˲'^Ƿ�a����y��筱�Wp!���s�Y�&݁���������#��#�n�)�*��vYDR�� �O�]d���j!�����ˎ���k���O?�[����f�t��^A"��H�!3G++����P���}��t�[֩~�\E�	�E��{�H� �%F�)'�{�����~N��	�܅��誅� ���h���Վ�����Ws�S�sZ�a�+
�^_%h2������/k�u�\V���&�z?c����d4�ֵk�u:�I��J�8�׏�Æ�� 3�w'���n�!�"��.{m�a�0�ED��\�ו�C��&#L`c�U�<�pla0A��S�y�D�E��++�{>��İ�yR�$����)��}���Tfaw�&���\�LgG;hgQ�?����>7�9��ua�.9P6q�esN�-��op�¬��47���9���L��IȤ�,�IYZ�MM
)i�y��E��GW�^�k��1�Y 3�.6V��_zz2pMP
�s�v�׿����������O�pv�Ȓ����J)�_��C��n�-�g�����[n�� ��K��R]� o�&/�kpsQ-<-�!�$����'O˛GNȫ�?#O~�q�|iVJ�1�}e��;Ͻ����}�:�u��Q5�ch��4p��l&��}ɹ��3�dY�̓#?T����ߑ?u��_j������q�::����5A�����[f��~緤B>sU�|�}�E�u�>�9Ci��p�_�>�qx���yT0��f&ݠÖ����ޝ��>(�n�,�l�(��,-�P����z^�۱�o���;3�뢮Ώm���LJ�\�.��a���1 `�����ª<��RR{��К&�	<y�Y�#f�,�{�;��y ����t��]�)0���� �4R*�~��������bAZ�9����Z��d�Y�F�L'���:W!����2o1s��ϹF9�a)4�*Z��w�����oțo��n߲�`�m�1�׷`�Q>��'�7t9�6���_��[���M�<�mq�g��\��j�}�Fiҽ��6���� �׼�ʏa�Q	���&��A���3gNӹ۱c���N�Ĕ� �"����\�)S�{]�u4.���� �x�����-d���ԯ��9�,��B��9�h����}M)뚶P�$�Lz�������
I.�@L9�5��9��W��$�����1E6��;1�,Ͻ����42��?b����c���"��|׺�s�k�R�� ��^���2�XKl��k�[�}�� |�B ��F�� ��#�aW����W�Ȣ�1q����W�pY��]Ƕ�:�TdF�IW���TGd�֑W^;$���mz\���V;p=�ݽ�2FQƚ�; �f:S���ۚ#���T���a�ʌ�0��i #+�}8=v��:1h.Ō��x��l�9ޕ�q���G�E1B��s�3&td�<3[��n���@,�����Gy���݈�1Y[[aG��H���92��hu@�Q��ԛ5^��C�2{9��w@Ő7JD���Q_�Q"i��F��`]�x�������K255!]47*� ��Sj,�ؾm�s��8��&2���j���S]��J��s��05͈��<8~�m�UG��+��(���$nw�E�щ�Ӂ�(+zsŲ� �4�t�&/h��M�ȇ�/l�M���Z��p����SP=��t��W���f�\��t�"C�1��I�%y��iy�{O��lI�����
%�f_id�wo֕W���:�v���Y�� �I��٠kc�$2V�k��Z��_S��G�5�l�8�%6>Z֓7eX��6���v�1*��kM�+ Nd�	�⠯WcZ_�S�R��N�����H�(�i�846-�8��v c��e�S�X7���?"ϼ��T�|��\9I���:�����	�|ۯ:�e��DbṴ1��Xo�n���w���:�c�(#()�#V-��k�R͕��Z�@6�@iH�� ��,fU!�s���$c#�����
���ۈ�n8ZIZ�3.C���(AkY���_��'e�:��!�!�� ��*����:���ګo��":������{�E̨uN>7��l9�&�'�u�n^�~�C�&�P������^` q���:>5�.-fbR��P�WǕ4ф�������੥�70s ��md�D�M�ɲڛ��qS�PP�356�f��g��'�mf�l�y<Z)��=0}�ɞG'������:
�8Æk��9>���ot�9}w��|���z�w<�jt�n��&ٷw�����#G��c�}\<���QC�I4�:�U���m���E����9������{ iXW[���	`���AП)~�m���!�*R�Ȝ������#�.�
2�{���;��A�_`ӏ~p���0�N�eyq��+�a�,BPtTU��Xv�&W������Y^?�l���D��ϖ���1��c/5�w���m�A$��e��3 ��2��>W�'��jO���p4� �V��K��_�7O��f����6�]97�r\PYv�We�1r�0�{M�6�9��o�d��2gZ港�-tt���Aş��đ��Ei; �#8�恞s�Z�-5�G|����))tS����N�^����D�x�2�LW7�Ē��S�$}�iy�S��7
�HL�2�B;Kƭ�Q&vY�&�T6x}˫+8߽g�L�O� �;���F<^ǴU�$�b�t�|����8p~������MXkj��L��r�ڑa#�B ;�u"}�k�Ny�ͽ��[�ꫯr1�#�91^����'B�h=oE���TX���>Ң��:H�� �i��q�������m�>�9h٣���<W��:�"�#{mYCk��S�lܲӈF����-�x����������	lx=���{e��\9�ōF���SW��q�`żacf,
�e�CCd.�B��;�����K�6s� FD�M. �uL�QZ���2pUC�r��yy�ɧ�}u+���MY�@�9t]�=,�O���<�\�e��"���Z�n�Mceu>t=�XwI+9�C�5�����K{�n]{m����6y������u4[��_���mN�k��&VntlJ7�1�븦��a��H�e�`4�!�
<#uVK("��ã҄���I-Yp��S\��7+��87%Q���06���i��I��)ih�꼬�F�A&]��Q;.�ƪcxp�#�]����=�ZoO3(��OA���#f�7� z�Ĩ<���r���n��r���(1k���2J�?����қ�e�G�#���\e�̧�+�F���k�2�S��}�'�HP�Ǟ��ϱ8:)�f�'_���{ef��LuI�V-mF�=$`˻��L��Ϻ�!� ��ñ���c�F������t�r���Ԣ�+��Kc�HG��w�'��Gp����i1��܆��_��)�Ϯ���z�^� ��ˤJbgk������y��妛�S���P��8{��7�	Bt��V��uP�`2��dǀL���ڙ�j8�(�zZ2�(n���A��I�QRVσ�k�kf�&�-p�n�_5ÝW]gq�9��;ഖ"���RX�`S��.��z��1��g��'��8�7n � s�8����(�xL��4�G��r��A�������sj�N�������%�
T��I�v�܋��.C0�('��w��['�J���NbjK��!/�3B��?{�]c���7�������0P�k	�L=i�T"���
L%v6�9���	�U�X���va&S�������e2Gڍ�!�)�t��R�>��w�t��`b�I��.Zx����/���'����Z�Λ�eE�
��6.�/�M|Z�A9dv��Ge�q5�sb3�`jQ���� ���� p�l��̍U���8�kp��2,V�x)�F�����ר���9ꡌ��2�����Fv����0H����;oс:v�����[��ah�@��!ՈL�u;w� x-g,>��Q~@F��{S>[����$�j�FG�g�%;��ڐ��2C����%|x�-�02�ث��ƙ�[Γ�v�8�N��I�3Oe㤈B�Y%띀4�p���9�tP.t�6�YCø�#�oj���ϫ�s�>�m'������E�DkJ 7�_!%�@�7b���Ұ��<��'�]u��������:����!��~���s��?gd� ���ejZ�+"�����`$K�@��X�-���M��*��9
Ҁ�sg��䫕&��8ȜD�ȑxL��d��15�An� �(�l���ID�]�7FFV�Jz5�ˌ?����Ğ1�Y���S1�VuB�D��LB���\�$C�
2�W�S��Mj��ؑK�\�Ǔ{�>�ՕA��pq��BIv��u��*���t>���x����q�0�$������=�RйH���J�zWƧ�r>�#�Dp�Rk`���i0��&	2Z����<�ތJ-c��=j5�s�;�1���s�a+�<q���8=yR�zoL�o�'Ude2���5� �ތ�x90|����È9�T�.*�p��	�?�$��֒zڢd<�ȱ��X���\+۷l��n����������t��i��L�A��~'e^��|i9wE�࣎�퍔�M��:�j42l��}�d�����nQ��?xB~��s����	����`��c�y��-���Q� ���Zq��ˆm�r������zM:p���)ug6�����5�����3p��k�-�v$,j����R�۷��l��h~�l��$�v��7�$��}�$�0H�^�k�n�[�Ѷт��n�ӁW{��+�a�f��8 a/��G��C&d�	t���EE�w����|��W��7I�:.qQ�:�J��D� �U���Wk$���k���s��-���l�q1_q��$cr�G.�([��m!�A�W���c�%�	�q��J����$�~ы�̐_}�mD鹩7R�#��ܬ���uˍ����@��j����o"�QMe����5nD�$�?�����QC�4�E<Tň����XC����eH�vD�q��v�0��ds��S�~�;�5�F"ӌRt��)�Bv$�[p!p� ow����-J�_���K_�"e�������g�Q��$����)�x�� ��hy����_"9�ejT滥���H!��ò�^?����O�8)s�f��w�L��k�L���R`4�vKC�FaϞ�$�UE�b9��|�4:� a���v��5���)x+,��Lgo̯�W�N"}�;�Q'�sƁ�d���@8�8�5���V����z)bM����p��v�t����n�5 ����o�#���s.KMK��t�ޢ��=x�����7nbf,�.<%}�n>�%���Gtm R��A��q��:#��Ʊ�%oXpl
)�IʬK���I�8��8(���S�r��oc�n.;U��$À, ��,C	��^��Z��Ӑ&���|����Ẻ8`x�/��L��"���ƙ-|�fl��C8>"�P�8A��n]:�%���@"<�]�,�ۈ�Wʠ��h�Z�u�KNDp��)K��x##)��������1�r��J����f����䊲i�F�7����d������BOk$%����9Ա���|C�ҏ��b�>�d��5u�Ll������&�+U9N����u���#r��4~�H��@6NN���K$��m�ƈ�GG�/������eiaN.m�&���%�S⳽����Ө7�%�#��L�:Ű9��eҬ�L��~���H�L�@=����8��3N^�r�p�oD�c�]=�09A���hm�CXʮ�8c�IX_�H�S1�+����V��XSa�`�Ǜ6QQ�I�I�f��
!��1���1X\\��;L\���&����*;�a���ܳ{��޽Gn��v٫N1eZm����� 0�ܮ�}�\v��8I���3�5T��^}]�1���@e���k*]�46!��W���ʒi=��@nvr�<���껇��6�"07`+���s	}u�g�U���F��w=�UFl}�$�ԢZ�k*N�M�'��������~���p6�W�Gy8���1Q�OLS�mL������h�Q�=R�E�flz%m���u�f&�"C8_��!��ַ]^Y��^z[�'g��Iul�eq��\��a!&v 9Pp!�)f�����lq� 0�Ih.���8.ӓS�|Bi)R��4'0��n�M��9�3nued��a�L�3d&�D�uoYi4�D�h�h]�py��-�f��g��I�Kl�hL������j��;҅�nm5!�gnߺE���o����E{��)�a!���Y]�(1�PWyaq�*&�gjP�Ӆ��(���ݔFų�G%0�R�`�2P1�B.E��hh���O�kbt\�)ɴ��)2��"{�eq��l�]dFO�8�x�@!����?	l���LA�c��V����r������i�� ,����B :��=��J8�h�*r�8���+�=�y��Z�u#� �
������5�Q����[fu���&��q�B������'$��'Ʊ;��I��g@����e�}���찖Ư�������w��a��Ѵ�[�9�H�� �K]�C���M�KX�h��W%�I���NC8��]�-�k����Y���_���,�����sO˷��_��Ȕ>]g��e��f���u&���sb�xd5�t�B��%s�,���
��1�p~�"4���f]ƪ ܫo�=�A�|e�V�{�щ˥:7�� ������u\����9�o��a�C=?:ȴ�+�rI�
��*5}�h�J4�i�Ҙ%v�Ex�[�iⰄF�c��C����V��H��g�m�a�b��Rt��l\�%
\�YMH���>w��溽R��S'�)�Z���X�w�J��m+n��B�Z�&�O�5]���;ddlXΞ=��
ʂ�:&�_@ե�Z%�k�:���3:6lc����h��~v8��/לԪ�[1���_Ķe2����a�&#�w����=�g��൱5���2���[ZX��w�-7��n;@}�_��_�#G�{���ˋK֌��|}m�������������J��1=���4j�:u�1g���-��c#��C�t�+���C8v(c?����@�}���B��s����t0� ��������'���7U���2U�>Oz)��t���{�	���`��`ỎG�!F��ɎW�<C�}~�Z�k��8Z�<�_!��/��Lu���B��#��k�ʏ�|_V҂4��Ձ��K��/L�ф�����_�a#��q�_�o�Nhq����g��Jm�UӰo=g���E̙�	S�&�d�66���G&'�lbQ�,�n3��(�u���'x�o��hӕ���*ؖ@d�����ӿ�[�����܂��YD��+�!�u�%�c�Y�8�:�A�tw�`��.$ =��K���F����]��b���D�Â��93̥9��sx��8��~fU�8B���ǈ��ҲX)��)�t{4y���izK����D^�_ ����e��/,+��|��,����u���N.��ёq:�x�&�&�����y��}��4�(Q�!���=�� ���q#
�Ռ�K��m4��躎eLdK�xǪ㲗q��8
�Lz`�Pv0�����Q�q�6T��ZD�F*rr��/� XU�f�(v��'�	PeW3:���wMm<��)��L�M�'3�6�!��:_�(�wy������#��ALמ����`��/=��z\�]�@��Vpl/]�#��Co��N��e)6�Ks�����Idiq������v���2����/�+�G战C	LmQ������ݳ_�޺A�N���Ƣ������aW#uнU�&���_��<w�E���:[mՋ�Z�p��dm���q}�k�a���X��aFsE��
d���G#Q�e(u �JV���|tfq�A?���9҆�9f�!Q�t��h�Vҍ+����SPl�xBvtT�Y�4�ܫe0�A��L�
ՖhH�N�Z�O���ܱ�z�Q���ʹ	�Il�~p����a(�k�%`Ü	Ւ���6ש0�թ��&����ծ��i��$�z#c�u-5�r��yY�����n���7�;4E�
eu�,�{�\T��'���+1~���3�������6�� z%P�^��u9�[F������B#�kv��~��M�J�-2p������(#������g���p��ۿ�����h�//I4��d�ꗯ�:��p1d�f@� )��� _��b��k(ʀl����l�s�-�8��<_GI׎��!P��g���W	&9�$�Z��t�n��4��ǜ���=����lƦ).֛ ���d'��Z�ih�N���Vy��y���ܒ����p�2$��.��0n6�*����b��4oi�}�������nr�}�;\R��Y��M�חk$�M���o -���\�\0���1���Ԧ�����VCg�Y��Õ��3D�Ha!�EL�>����o�׿��04E"�0*� H��8�8Y(�v��kH��Y�7 dM�@F'
���:5��ȣ�$�kE�EDҲ�P� ^
/�����ҰI:ܜ׬<���GI�Ge� ��� �%}]�������ǎ�1��;"9"վ�n�p/\�(���,-��T:MeD��Ƙ��N���D����u˖��IJ=ı2��2���e+=��pP[����ý�v�uf3����
��԰Q90nLO%9���~�8���>+�^�=����B��[�7 ���I	�.<s����AY��]��E'I���(�#C�NLdch`���	���.`� �k�C�sZ��:z\���I��|ɴm�#j�F��$��#� qM��;)���$o�u����$7���!���ȳ_�K���6�m�4\��tC��R Ӱ�NR޺�ѽ�^��w샹 pR�ևw5B(�.]��ZS��D��l��?�qy����X A;8�f���6�'K�u���g���\�:�>���u�\��z�!�.��d%�K����/'N�����<1����r�޽�������^kj ��H��|�l�y�Q2e�X0ُ�\?~��=ʷ�8�t�:G����&�~^��0^��֗�4h�sU�Y7��.�ʝ��;�ݒ��̰����s�^l�	�6(k�ɥ֔��r�&V�z�x�EbT����-���/�N_�3���yLL]�M8���X����S]�d�22� դ�b
+t���VW���@�YǤ���+/�(k{���۷I[�{Y����e�2,�\��q����`�hvB��5st�ȗC?:0�F�ޞ�iM�w���LW:d5����]�p���ik�i����?��a�Ѵ
5��DP�!�H.E�_#���1Q.K��y��g!�%�895�}d�����`��]�7��G�f���^��s���:�>n<�]d���e�|菘��w���r�э��xȱ�rM����T?g̢��9��"p��(�L� ��~&��$_�K5y���b�-��Q2Z�y�N*!�`��f�������$����j[�@EǗ�C@�\��t�)AQ�3�����&���K���uz�K<�2sA��IT��$Z�o,�����b�e�H��A�!btJ/X���Am�AL 	>$� �!�чO�%�����"�8����.�4���ڀd%$�y�^@\2F�s���Ffx�b���T��NC��`+ygRp��9�t]A�J7�,�0CV�ۦ�I}�բT(,�il4Z��4�Ƭi'��������2�4���4�{�sG��F�\(?���2��FpԻa�����'*x�e��Q�V	��F*����'=��>_(�ߔj$�:���D�O�t}?�Äq���^\����d�ɼ�g�ٿ�WP���	�ܵ��Q���H�&��BR�yY?���iE�J$�����HD\o� ���.3"�ht�5�J�N"�����SraQ�0h�F9vS� ʣ)Ŀaϑ�JQ��ϏW��k�eM$]:Ǡ�)�����r���j�'Hd�����<��뤥A9�֛vɽw��rE��kRW�wH�9s>1�x����ש�����	�usZ���܀�jE�����BQ)��'�A��*t�i,S��t��?�������*_���J�������ߑ��-$�n��}�=w��kvj 2.�V�dX֎+�v�/+���$�����M�L\fN�-4Ik4�膴I7�mSc�&YY9)�%
) ?��t:O[�>��¾�W"�������9q?k������Bʩ2�0��S/j0te��2��R�-�I`C�0����+-����Y�u�?J����Sú��9AǮ3Ց/U�.��{��s�uy��#���n�L�M3S�n�Zcw�rc.�[���G�5"p�2�^�G��sF�K�؃}0�Ő�ʲ�(9��漀���� AHu���Zl���$m�A���6"���j*D������:ܝ����Xec�0;�8�Pd(_�O�H�� �{�ڻ9'�J�9G%��8q�|�q��@���]��	�3�^u��:�C�'4��߀����.�YуI\p]ld�2'�V�4'1eu	A�R@�4\it���w�1Q�K���^**z�ı
�\���%��go�q�|㠃�1�z�{�0���2��6(r8�������Q}+z��F����D�>K/#Վ�`5�H_��n���zl��Y��b�g��d�H�N�E꘬�4��R���O�<$�km�U5�c�7�%ЅA,: `n�ܨ}5�ԏ{�c�L_��z�B�E�)��-�*R�o��HM�%�%p��Wb�����D�"D50ڑ+#�F$C���'J���C1�ɘ]�օb$��`�< 㪎9(W�9Ä@y��EE}@�p�l2%N�2!��겍�sia��w _�5j ��`j|PR�7�u��L�+F�&�����M��6�P�N4=�x�bGC�N`F��8���h1��'�F��� 3���j��v=	;꽁��
d��
���Y�rhJ+�оM���ν��.0T�@ ��8;�,'%�tSN�V�%�>#]8���҉B�l�XV��-�\Zk�%DM��y�Կ��O��HŸݠH�:'+$Y��H���'���3���q�Д&�c4��H.uu�|쵷�S,ȿ��gdttD���c���:@"9鼞��j"��5Yl�9��1'Ҫ5h(ӥ��id��L������� �hN+� h�4Տ����Y�����:o��Fy�K_��y�{RPG���\�]� ��I[��?ղ�k����nj%���O�6��S��y:lc�HX�qx-���_6M����(�{%���ߗ�/S�s�AZ)'?z�Yf
C��X=���A�:�݅TƆ��{u� �jG�n'�5 4���a��w��5�}��m�k���G���:Ӌ<��3�j��g���ZS�٠d��r�֠۠I�ԗy��p���s�&�����;G;�o�
-3�nR�剗^����O|B6�-��U�ڦf�O3i���d/�("���~o�*Rp�Ѐ�֑��T�ȐN���/��Oh�-�m;T��7�c�Ve�~L��B�@��EB�y��(�I�� *��
�����^5źKT�5Y�1�Sb?��Ob�K�e�@Dι�cU�X�֜<�s����ܟfH��N�-��	(�ਯ�Lu�d�����zϹ��-8��/\(k�.p�|v!gU+\��A��"�O�^��;iı���x^�>G��]��dp}`o"�$@��!^s�7��aG�LaCK��t>��I��l�3��̄�;�{�����wQ�%�H-��8ܛeV��G�xF�<yV
�R#S�U�]�����]�d]d��֎d��)	=UN��g�Խ�2�!�ם/�F��hAdc�����ϖ�8GJ�.6����L�v�F��8D�4���+uao��U1�9H{;XW�H�!����Q�Ҍ�sG6/,��15������ÿt�̌W)|�F&z}͕�M��!{�}<dW��L��`���%����1NI+5��E��k���;�\\���31	��#݃���ĺ�\��D�rg�5���!*���9�͇h�vn�jvTEA�GNc�(n8X
�F��fs��Yڨ� �p����}�z����.���p�r�GYF 	\��z}�_�Ys1������Z�J3���$��i|F�e����5u[+�M$�[�<e�����s k��c�u@���Z7aS�reLJ����1�y�cj��o����jA�I���W>����X���������&�9�`�@�uc�c���ߔ��U����J,��7αy�V�x9��7R�ӓd"�Pg&�O_�:FA��;����0����pL����b:�a)���r��)�a�4������l�����R_�,�ڂxM׃�e(*Ш5VW<�e>LB�*Gҷ����V�B�v����l����n�Y��E��]�{������a������4�vfZ(q�#�88@�i��J�~P�R����o���@p=�{�6������[�YIM��s=+(Y�o�����OH��u��k�J�t]�m�����s=q]ͺ��|��Q|�q��f����MpPX� J>5��q�h��X�U]bg_ll���i��yf���ge�K �(��5�?�a*��F�NK.\�$g�]������(ռ5�S��N:*%�����  �lg�JT����ny5�.�Y Gj��2q�f�n����7ʜ��?�w)��q��J�v�Qoy�����%i"b�g��&c�6a�s>f�������A�x����c�g[%�|^e�䌱� k	b�\h�i�����,6/��&���._��?���{R��.+f��I�ti?e����e���,�u�]�#·q�E��q�SK��?��Uy��!./�\a	��K���8��8Ft�bi��l-�Z��F_��c�٦Ƒ�l�� gZ�tq�uO���AL�"۞a�y|b����5�k�Fv��q	��ʧ�C�����x��zB,D>4�5,���>�d�a�ePb��IOL�~�"ʵ�զ̶g����i
��-p���"�-%~�vB������@���t,O��	���qs?�(�݆�L3���I��tH�l�_�!��o����\��a�3�?yW�M��t�}�~\	���\���}ê���x��O$�Ǥ� v&�h�U<���6��L�����x&tf�e��\)�4H&b+��U��<l��t����R�/5ǘt#��[����f��{ei�8&Ò���֑����9��&��K���ݴi�9:h�p����͡o
|W+U��/'Y�+�f
E��7��e��)y�����lݴ���Nb�'`n�WT�xG罹�3RE��Ij�@7�r�6L���t���������r�q������5;wI�]8'��`K����C�$��IJ��\���7���ɵ�.�i����u��2��{Eo}��j�z3I����������/�����^����}_���-;$7<*�-/|M�ݲLML���y��J_�0p�c��˔�|��ɸ�y	P�?$D ��u͞���7�{OF���@���K��'���ݳW�.��&C=풾�����U;R� �����l��fe�i����=�3�/W
_gڰ�*V>�A��8"����Vw$��)3c#d� t'̻n[k �Y���IBGh�U96���:�:ǉk��f=5=!#�����FruaQj�5���� lX��H�B���ʼ\�kF��	�3��kA��y$�� 	U7�C�.O�o.��sh�6��,����Ճ����:�0t,��y�i��Y��nb|�k\C�ZIܢ�Zwn�%v���[?+�sQ>~��G���E�Û.���>��;�����r����f��h;�2����8��R8�:��mG����p]V��U���䴜_Z�o��?�k��i�1���6��+��[�U���Y��ܕgp��>ۺ�[�����̞?v���'r?##��j��KE=�Y�ښ:��&�1�j�6l�J^!�	=�Ч� o��=����9!'Tإ�t�� ��M��C������r��)W����e`���ojy=L��������I�p�w�Y׫F�3�)���hU��#l���I@��%�Ԛ{�H�#;C��С V�tF(Efj�l�������0y�\/�H�hdl��3�>kh�cb�� HO�Y�Ak	��A��u���,+=��Ƣ_]7�0�ո:��M.���D���2s�J��_�k@g]��`��S�� �X������.�aK�.0B�2���Gd`ч��XƱ/��cg{۸�RqrNu@H!��P�izZ7��_���\��:9#�j2�ߛͮ�Z8Z��g��w�y�0yW?	3�Z��~��#pY��G�.���0�'j�2�kzI7��=�#�a�ցY��f�us�JutLF6�Ȃn��VS�:�K������P�q"3�_��8�a��
Vuȇ��uݡ���d@�M�PJ�畣��߱C����ٲ}�9vN�~�0;9��h]��j�+�ң_	�����'���_z�A*>��<��=i��rf��ML�s�N����+8�p�M�#��u��\������di_f���>��$��#���l����+o���"�=��Q\�,��B�\�}�@aI7��Ԛ+|��.�LG�sMz�q��2H�+߯Y����F��b7�Ss�*%���{kA�=v���O��q�>�Q�f��
ʅ�����,Es�A`H�Fů��c�֖IGCV��(tEo޴Qr���D����z�T9xnP�0��H���\�]�Օٵ}�lۼ��jU@a*�0��{�a �i�6t"��OVY�;|�!1���Y�4/��zx{���v;�I$nEI�jϻ�Ƭ�>,C�I	��ณݡ�8&ͩ�\�a����O�A��`�P��6w?!b��e����?�B"��s0�Rl�����O��w���Ș\^^�Ǟ�����5-���(�����N��J�u5p\��T�oֿ�����p���>�A�øR���<�w �Zwt���������T�Z�%�OI�k�*JR�RWc��tmMf&��7$K��R�|Q*2%I�(5<�|Q�d�f��,d�$��L#Qā�CxsA�]�J'(�b��l��HY�����*��^����喝4�����%�Q[�yl��)h �0�٥N��jIf�$f�J�=Gל:��vS�MK�\��pk�T1�W7���v��Y��+�#M�
��È:�-uH��s�[>f b�I?��v�	�tq�wޕX3R^t��� �C��-\g�t'9��u�y����&�q��k���#�(X��」�y����KR[��S�����?) �h�I\9��?�:�����Ȑ�/-��Y�E�'})���Bm�<�(
����v���41���e�mu�5 98l�_&�H@xf�S{V��I�l�zr}��R���8�Jjpѧ+3��ʣ?zFy�)Y��P��*�a)�5�R�9���\�6ֽ�	��{��$�ʞ�ͯ/I�
�W"�Z���y�����3�mfJ��8FbdPߌ��K����-�Ȇa)���B�Y�
89�k�T� z�&��d1�ƴLH�e80KCR�N-x�rE+��Y������\�Ŷ}��=w�+S��Κu�c�+�'o���|�\�]>���?�gr\8��<`�����-αv����S�R�߁׳Y����2����_n�{:D��ǿ������=c-;�,�}ι9��*�bE��%*R�ҴZ�Qݶ�q ���/cx ������<��餙V�[-5)R�H�s*��Y����7�s��Z��ν�UIbw�@%V�p�����^��[R[="=h�aGV�l�wt��Ԇ�r�����8�N��#���ϟ7T��꤯te�������n�dS����!i�|�R�����&�,i0��$`8��V7����ت����J�[��_L��F��jk;8$�4X�$���Ժ�"�o�"oC(aTa?(U啷�I著��?�~���S� }R7�?U���-�:�`�+�]'�ɴ:�t`%t�vc8z)M�?�ys�9 �G�qp�QYj�������@������r�ѣ�;�ҽ��Jo�;$ERJn�nI�wJ(J�I\�%���	~�I��aF�N:���>�m�A�7��0�M.Hr��y�~F��<X ��'��g	j�9���	���
̫x���/Ԇ��l->3����d�s'Y`����_��?f ���>ZR���_ϻ��Xs�qEgd��
K��C��mgí#ݨ6��4��k�yk�%��?~U�4Y�j#���E��^3`�(��Io�=��j�{�l-�{��N����Y��#�Ͷ=�5�Cf��̚q������|'�ǃ�y(�9�kj���b�am#G��1�;Pó�l�|���h�pH"��)��d����C=��g�t�3�Oev��Ts��������\%/�v��^�չ�ij6����ⱀh��V�+��o�J~��_Sz}	]��;o� st����kK�ul������=����vIo`��9���{j�77��4�{���Jނ����2 ,��f�]`�1<~:-p����xIB�f��K
MK�㪡�����o�&zHK����).0�㚐��F�����áVC��nl��N�})�SfIHA���E~܅	y�ԁ�sPn/�3�v41S"oH �kU��\�5��ǐ�dhT7xOr����M�v��5"�j����g������e
5:A�(�r���2�H�}ڝ7[s����IO��f����h�z�$�q�ƚ�Mt?}�}�����h7�6�g�?+�y�q�\{��8�X�1�	��0�C��	+BH�0�����Dx�k\S���u}jK+2�~!	5糰ojU�i��QYFJ"u�5�o�-BE���̭.K}I�QY������8ߐm]��z���zoo�;�r�I�!��� ��?���;_�Gp��s�Ƚ+j�������5�l��Uf(���Dܜ#���^����v.���D���4��D}��KwcW���o�u���slݣ���h�rU���'�=���?z��Xj��F��I�a_�IF�Z#3���^1t��3�⯾,pI��z���Y[���k��ܺ�(�BD"*�9���<Xf&�H�XZ��[p�
��>'��\�kG�ee~�������K��B����4R?��n�����e�O坧NIs�!*���a�Q�/�Qt�^%_�s�Jf�9�F8�/-g�
yK��E
����~`o��q��u�#����� wr�1�	�7�� �]7kO�y�:ٙ�>�Q�O���i0���3�������(t1<��|i�BX+��������}�bGCNk�R/%$�PbtHB���J�?W������rv�X�d�DN_D2F���e��ۡ�~�_\��?�������q ��8
�<����`g��rzP�/�ҏS�	��*B�1"�L��\��	(�e�,oH+':�$L2t�:g���i,���q�&��&�q���,^q��UtQ�H{o O����:�"�w�C*��~�;
@�bc��47E�&��$:�������X9l�R��!�3;��ʉ��la�Z)TX�I�|�l�jv��8�O����Su%˘H �"� Z�$�;��A���w����wRj#P`�̟��Ȩ���9kD�Bl��m��
�A��]����Ȕ
l�=%� ��vYf6�u����7r��`�4�z�TEqUg8�R�79���w�\�\axB�q�&�QULl �dF��8w�5��L?�˻�j	�F{����0Q�;%���ȿ��o�P�
�օ������x>8�{�됒�`2q�(�9\�=}`�}�tN J F#/���]�:.��J�&w?"�VW��s兗ߐ�nK�Cdj|�����JP�
5y\i4�Z��ںc�I;Ɩ��ӂ������h�U-�8/g.^�?��_�ɹy�3�c�KsU7d���B���W���u�[^��?�D"�h���ؿ���Ž�9xg���ԭ�5����?���Ӳ��n|Mj��z֫��v5��6�t�C��e�Y�E)�-C+�Mn�;8�'��M���4A`�ΐr�#����~P�US�t6����y�IQ�.����C٘���@m���`�}�-��GDٿ�q������ݱ3D�K�_K�q�+�z�����g�}���WAX^v�;z_?������7�#�����Gn;~�R|�!��P�s�O�ɬ`��c:1�؈8�����siu�:�r��4y*�˯�v�"e0��#������Ʋ��'��Z;qdEN�X�����		��Oa_F}>���9�X1�F4%P�7�<����홤o+����z�܂�/�(�h��嘃S�7�9{��=��o�B�⫧lG��9����D*^#{zC��
{�)$�m'=:*�,�����&��&��K��CL���VչM����{\^T�j�����M���7��a����ʹ��J�$�
;lms?AF��h�fy�s�uŅM0�gى1�cJ4��Ā����浫��m�o�I�ޔf�&�`����_䬍y��L7`�F`�f�'چb&����U�rjD�c?yV�����-�q_n$��4<Pd��̅V)����n��8^=�7I�����A��]�cB�Toh�b�sb)�}�Y��q}Py0pß���|��`hu�P1�t	�����J�e�౅�J��ϓ��l2	I+�������TVg[���2��r��q�/(��z��k;�d��؞!��H��(����7!'g+Q�.&��_�Dܠ,��p@������a $7�C�&���vk۵����D-�0���j���ȼ7�a�%�?*��!	]�:��|♗�/��}i���1�j��� v�?o��94�=O�w�gZ7�:�ɾL;�4�ߞ����1��s�^�V�#���R·�ُ}P�ޞ�UJ����쵇�&d_������H{ؕR�F��!9�bzЪ+�zH�D_����m=;%�_9*��g�(�X�X��\	�^C������^��/�%��]��ms@��:/+���J��{���E���u�#@������|0@�VjْwD�p�a+K�mw���}�|��58����q/�ﵽ�b�8F����~�����g��l��L3М��p0u|����4q�Y �0�(���a�o��1=+���i��qmC�Ce�h%�W�W�W��t����H*]��v��*8�\Z�/��5������W�������f�(1�4tu�c[_�TQ��,�]'���O;9!s�1�70���d`[��vew�#_���j���!S��t$/���D?^y`�����aga��B�ٿ���	�����}ם��k:�L`*Ś��ؘ3`o�/Fݾ�m����	�i��5`\U�P� U�|Ā+ү-Y��X��sC-h�����*\I��������N ��`~��� ��� !(���߻ٳ�e״���o�2��܈qtW5�]��6o���b���?��v I����L���{��p�	�Xx��kץ�h���t�C,�4��~M�V?����7�'?{V^8{N����w����CGq&�k�K�*s��~��)����L}�t�41.{Mb���5KB�Șfgv:��r(�z\�#�67	��J2��S�X\:j��0�u)�+t��^M c�O�,���k@���m�fZn�f P[5�)r���d(��#��X���-���=�_���G�zO�rC�rDz���!����$��s���,X����ڄO�=0��{��Z%�zc~���9dVc�8�q2u�QP����RV�Bг���@�֬���)�8�u ��z� KSag�Z0��l�[�&��,T7slk�|-��f�*ny.���#a�g�%�T����@cvN3,����vMz݁�#����%��=A,�uDFMk\V5e\b��F��a�+����EY@m:���ϰ3��=�}?qUd��w�*[0����VXm���g�[>|O����p�����J��&���1y�ɟ�^��LZ#@5�T�����{�L��e��Y�qm=� ��q/�/�?HX�T�f��B%�w65�}�rp��.�sԤH�I�g?�y�;��g/�_����ճ|��H�S$a��FC�sN�g��kMMZt���'��ST��c7`�Ж�sA/�9�(��\��_ҠsA`@��\��5p�}2����J�Hv�n�ƾ��3�(�@�~
AY_��&%���O&�C�])"V��z�d�����8)���e���W~xT������u�4�EXJ�ߋ{��sD�L��mL��x�`_�~E�9�uн[���o�I}�J��74q�棏����dE�ߑ�Ey�;V����2��S�{����6��{X��xI���s֊��MRO�فd� �H�~�m2%.&X�F^�x�5��.4��$ðe��d!`��3��<)m��\�[e%��3��������4������X*�L�0䞲�=X�0�g��YXZ������l�*"Y2�X/�؊��E�g����[��ݑ�����M���X]�!��+����Ʌ��[O��ʲ4�G�77��.Vʚ�|O�'N��	�v��^�'C>�\����{J�b��r>�7'�ϗJ���O5[fk3r���kZiE�of�1�t�A�,<2
*�V;^�z4C��c2�)4�����֑򼓾Ce��$� GW�h`JE�S׵��[*r`3#��߫�s耪�t=�6Oh�@�
t|��=��@��"���sO��y�ŗ9kP_=.{��T� $p�3�ÌP{_yC��`�����9KwN�?j_ڊ8`f}��>+�D�`|����g�:��{θ�k�s9��I�1�m՘�*O�
lM����BŰ��0�B�p#Zj%}u�ˈR3P�?h�\%�WE�7��c���if�Q����¡c��ِ?��o������#u���=bQ08b��+�P���S�9�&E�+9 ݃EL��ല�j\ַ6In��#�A�Pt��FZ4R
O-5)�8ӨD���k$����=^����$���z<	��6�h�i�V-���:�A�L��&]e�K8ް��n���y�H�"Ǒe��O4Z�6���<$.�i���{ܐ������Q3�M�4\~(m�G�̆�����񹁆E�?2���)�e�#O�؀�o�`�
%Q��Ac�J
�|��6�}0=y4.�^@�
��|�����ץ��$�IC��%��nl�϶�g������}5����h����;ۮ����fX��9��|�o��s5���}ש��_����KM�����&'��e��ç�Kk���M?'��t/�t=���ĳ�A&�@� V"�SV�2q���4�����U۳�AnM���n[�|�����&꜏�9��!�������OȖ�d��6$ĴK�Ԍ-�A`N�F��+�G����f{�����mӍjU��.�4irz�ѐ\��63�;���X?E�'e�B�p�R#.t}����fk��tg<B�:��{��&��驳�]�W^?'_��O���I4Cj x�ʚt5 <��_g�m(=��s��~��@h��7�2PG�
�����!\	)�
�v��8Cd�\ ��y�*���{�-�9�C��YDtz��P��UC]�N{ ��O��k���,
4�M	&}����L�[d����Н� ל�0��G#���sBV���00�j�0���`���N��i�AŢ�"Ɠ�l��e祗!$��<!'N����&?{1
\��R!�MG��Ï��(��́���K�����ә��<����Y˰���|u�_��Z��PG��=������~�a�O�D�����E�����/��$�6
�\�m��i��ǡS����#8q;���� ��8�� S��4�(�� �E���(���D�r��k�s�Kr�ں|�'��W���b�C`���/t�Ù���8��Ac;����7��M���b��0;�<ˮ����Iac�6�Q��_�����vm�) �T��L�k�J�p(h�bhC��o4H�!>Lh�&������	�_��n6��/�O@� �Hj�Չ�,�B�1_f���S?���u��J$�� 8��={L�@1&'��*q��׋Ր$��F���X��!M�e��C��C��J����<X�5T_`DH"=1�"*�Ȉ���2
bBi��9�M'��}�� �Fp�gK�$�&�������Ĉ;#��*&M�5A��RG�[�>�;�sS�0�k�j@&��iw{p3��� B�nө�@���t��%2�o8iz�(Y���c�s�k"��g4;!%'��	,ib�s���D��we��¹�귾%�<�s	sR]X��vO?Z�ؼ ��9��Fx��mB ^>�Mا�[�Yِ��]�$�5	�ȡ���U��T�׮oJ3ʙgu:���'�q'���_��������$����jp�{��74�qTCM�d��۠DB�z��Aa������x�;sg奟?��mAʥ@����GK����9�����^[�*Q<"�.,����	��;[��p��q��03�!Fhq�EUm�uOue������\�j= �Cyb�ݑ��ݦ�9T�X�1�%؎�xh�"��l����)d����b<�AM�ȝ)���PmL��h�Q�@eN�n���W�dTG��,ȹ'rf}S���z舜;����w�%{þ��S��ۏh��}V�ހP��YJ�nl�~�Є	(�FDv�
0�\�d:E�ֺd���n��Z�pƳH��4�
9�'*`C�KI$�]k}�G��:=���I9�Ԕ�fM�w���V ��5C'�N���g8XhR��nO��8=DMN�jb�0�� ���NW}�Dv��Y���6e�Y�D4��~J&��@.��kR�+�rUN_�S��χ��E��)Q\��ݵ�([�h�2$E����@���:ɱ+X�,g����E4Z�
b0�m���`��~�Te��D�"j	6�Yr0����l���"�7��;��`����{?���g��'��4�s�/���ݖlnoK�ߕ�&�� v����$�Z	7�GVm��x�_~U�����Vg �ʼ�ii �`�ClH2���~|��|�{րY� W�����a�	q
���#��: ��kE��"�d����x.�tQӪ��Vq�Ǒs�"� �*`���G&>�V�G�K^�_�A���n�Z�iE�H '�����v�˄�'RM!��.�WC�-�rcQ3���D~��hD���O�{-��Ñ�{��Ga5�v$@𡓠C�(.�<]Dj�r�J1xB_��"�Kc���ЄҬ�y�K��=�T��j�NKBF�$*��1<�Bޣ:Z3X�~�:��abr�8l�PO{?���o��g�O�-�;|��7��0g��9��������=��������!�0�GЊ�n�?V#i4[ܬ@��z%ޗ�P�[��V�f/@&��7<|�@�U��j�&��Ij��������;��e�P����9�j�`���)�1 ΅��nȿ��_��7d��	���\�kS�΀�V�p�X�!��gb�6���8����dqe�ϣ�ϥ����:�xo]�9"k���B�*�������Jqq^@Ѳ�{]�����Ƨ�iw�غ�G}�C��f���ߩ�q�ڠ�`:���n�/��g%|H��W��o����%�_ML�&�,��g>+_��/s�������.�F�_q����wVi��"������
���zk튼s�6&:Ks���B[s4�� �|�"�����h�i��B�����I@ۑ�8�Z��tl�,��	�`���s�Z�F��(�-B��`a~��I��]�����$��mp:h�RQ{���:�W�]���K{0&�?��+*�i��M`k#rlN�}��ސJ	�b�0\�����H��iE#�6��dL�8\��ٳI]�U#쟍�=�_Z$wj½&l�]�"��N����d�Y��E@�6ض(���`46I#�L+�>b1t:H(���@Ɣ5�I0 ��7�D��o�n1�\\^���E�h��®��U�y9w�\�|In;q��J+L��/�9��;B"4�� &+_I@��}<�Ja��x���RY(�(ia8(1l:+��CÚ���rF��3�b�����C|5�������l;T2zv-ofgh��n�����	X��D=��L��S�^����;DL/�Wjm��&N&�2i ׈`Y>]葉�S����2�-ñᄣJ]���S�=�y�JsI�H��?K>�4K3�)��K�8��n\ }!���6�틋fm���1�����X���nCb�Ù�����'�L���#�(�r�!8�9�����0p�"P>`��!JV�M�d�����l�|Y� b�帪68'�ĂK��o�L����E̩b�l~���M��vp	9k3 ��.����T@k��喔v���c+��|K7#��9/*�`��F ���G�v��&��W��=@u�G�<L0�(�#�������ŏ��������������U��c�.d8f��R�u,Z���M5�\#��UKP�(1��@j����yS��G��ho�pq�.������]�%˻2=���9y��0���x`��8{�=������>������f�0��jf������:�	B8`�ir�*D�8̑U��x�����q֊��T,�a�eb��>��D`C#��l��i��?u���y�x�ݭ.�گ��se�A��`F��X���X`��?!?匼��-���R���Kž�������^ĉLϽ��Ł,� ��g��Y��)b2cU;���K�` Pg��䢪�5u�G7�����u�<t�}�NT�hո�5����E�����Jd�A*TOD��l�@����F��#7#��v��g�����_��������	Y-O�Љ����.����_Y���c�����}�Sr��]�|�"[�R�=����^�`0-����I�Ե&��"^N0���Lm��#��:�Mݿ��;+��؃2�6$��`��vG� ��J�Hy�6�u��QF���vm��+��N�r���Q[h�~�pXC�1���i���ۉ{�l���Y�B"���[c�)|��ssR�5mmi@X%>yx}Kʣ��v.�<%��
�^�v���S��[W�������Ҡ�X�t0�J���W�ޑD��R�������+}�h��ɤ���%�BC�r�61�7l`b�u\�<ǎ�;����e�HS�jcY����n����?�WΞ������-�+����.q�pLj�����(r����Z-��K���?��$��a;֠��χ�1�M\���?�Tm#������=�@�U�����Xӗ�i�um[V�eQ�S�R��X`m꽽}4�q���v9��Ӛ �l��ɸ�]t�8ăna�Jw��-faMn���<G^%%�AO_c`�8��$���0�z�OnP6K�ץ�8�$%�2ř���T�Y`ղ`4tT.�P�{%rxV��ѥ@����v�
�xk���h_�!|MK�G�`M�s	�N��A����c�K�LJ9���t//iru�בo|�;���ϩm�HRiH{�cr�8!u!^�8�O�����L�;���8p��d��$c]g������P\'f���*�ʿN��$F��F�ge���k�l�XmS0�G��o^�-H<�!'�� �����#S�@�2�%�R���<d��;=݁юnpȵ���ȍ����
#+ nA��3��8b1Q��fc���ǟ}�����r��e�Z�Y'��&0kf�t��d0"��`���ͥ����C&���p�Ӿ|�����mNʦ&l�j#.k1��aq�)O3D-Q�̒@cp�65�M'�0$�/�F孪��E<@�J�\{7y���Rks���H��=ƃ���yss��ژ�L1���N���"�np�=��D5�W>�ء�g��UT���
��$pr��K�od@h�`?z�3�u;��oC��'� �ɰ�'��)��G*l`�/1x�'�Z���$}}�sk���O�T�|�U�b�UI��Ďo���/��}.S��������[2�-����ֵ������u�;�< w>.��1H�;�m9��9��ȥ�]y�g��n_�Z�AUtCf-3��*١c{�!��L��k����E���1)���ݺ&k�o�{�;����?��Ύ\�vM�SRj����D�_m���5�M&���|��F�eg{zfnvY�����t?(�ض�\�z��IQ���g_����rM���0�g�ǌ��}���"'���P�vkO��l�D�fd ^���w��x^� ]��t}���MB��\��b��C�O~����w4X�{<��(��nVO�}C6�9���ru�'��\:mL�/H�6����3m�لz�6���N�P���V���y.�8���ё�#`LS5E�o��aJ�֝N��8��+��S��i�x��~��ξ)���T>��3�� U^Z���B!��T7B��&��uX���S�^�8?6��+~���pH*p;(�=�"�+���i��eo�š'�w��� ?R,��Y����'�ꁛ�Vٺ�yLr6�G
wF����/�������禔���.�Ó#i� �8[���nu{lK'F��'��;��͎�ޣr�t��4Y�/�@��d��-�F�q�"��掭�0� ��y�1�6e)_t����X�3�������h�#��ڕu[C��$�O�uX&c<����V�F��J|�A���޼$�}�9y��9I�M(B��B�!<��k�f|���N��h������'NihAb 7����Ef�$������L(8o+���H�,7��]0��D�j��bGc��3~�Jß `-� ��x`�fC6�zF�E�Ƌh�%�8�R�Yې�L�|p)f�$�6�=�1r ��E�7Tf�2��'��:�q_^|�u��Z���w����S�`��Q�qM�ʒ���9�0+�cf#��ko��=���D�2�s2)4E�BTfp�nu��G��]g�n|L���*��Y����� :�duB:�H���=7ƀ�����F>�NF2N��oѐX0��m�uh��@��k�X�~����NL��41)<T%ձ�^2H���p&���";��a�P	����B�ќx#���A�	�!9Y��z��ޫ�X���L"2W�xd=7f�ߓ1�C]j�����A'�<d�BU~����|[6�ԙ��j��]}l��r(*��@-f#V,�[v�P&3�ӿ�5�*��b���ț�X׆砤aN�G�y�|��{��¢]]f�jW�w50~��K�څ758�=��E���i�ٶ�]�&��)�)tU;K }��Ҧ.�,aڰ�%��g��:����@
��>�P����8,+���[n��ݖl�4(V���m����5y�ʚ�v��t.^Ѥ����)w�\�9q�4��a��z��t��}rZ�Hj�_� k��2�zT֯^�0,w�x��mwH}aA
�y�Һ���)׺��qA�R��fO��u��!�9��U�,(@evVw����X�� ,���yV���c�����K�^���P��oJ~n^~��e�>��`].mn��EjM��,��c� r�|b�$�'`1��wL��T'���Z�@��������.+�:�� *��\B���y��q��\ފ��'R�����ݑ�Ɔ�w7�O^y]�͎|���k��23bMCMF0ąT n�"��&U��Z� NH-uӖ�@�s��0��FC���Ґ�(�zd1d�4踨�5RU�Z-KI�QB�ј�t�N�;l���"!1;�6�]�ٔ��C�2Q��ڐ��٨�UgA(>����{��a�.�s�鬯���T_���N"��ڜζ�ca��Rb4ݦ���9q��n��s�B&�U�4��GBEm����&O��T"Zz�>[��$�y�fn��E7��ݹ}��x���A�V�ͩ�������'��G�~F޸�.�����q�aD�1��z�H�Nf>o�!np� ���O5L��Ѝ97�e/&��?�P$�,f~f�>{$���kU{\=x��P1ß:F���*���`r�|)w�{�&8]�Ŝ���֕%����l�u���ɾ�7�����!2�@\P�j���o����bk�Vbӟ��Ѣ�\c�G$J��ߡ���r�[oɷ}Lx�}��ORә#�B�d�vl�#��Q��0��A��2�9* 7-��4u���c(��(Ż�FUKng�E��k�[[�J1����p ��tznϸ�\{2uk.�g'n�XkYЪ�aY~HY#�g�XLP+�Tv/���� ��禛�L8�҄+��Y�1�ơfU�\s����Ć8����@�%ʱ������1�tM۳�\��+�X)�X�'u�.>��R��G�M���ʕ��:���q��5ARm��}R��؏��NO�xo�L��(][�P$�q�?F�f�fVMc X�.�p���|�����&�/�������`���My�����<#ԀF��!��0e�ԑ�����7ź���{O��p`����f]��]�?��?�/}�r�JMj����W՟=w�����&�d�{�ӯˣ?{V^�tI�G�h<Vd;���%p�l2W&S\+� a��l�_Ǣ�p��jr���� <"����k9t�&��|y(Tc9??�kQ�3��ʟ}����kgd��q��5Ɔоn��\��xJ�%��Z�x�R�s�w8T0qF�<�p�;��$w=&�R�����?�/dS�ŋ�e>W��GV�1���Ӓ�_{�vqu��@ʹ���-	4��=Z��#�Y��t���(R���D���q�<�ԧ�%�~2l��S\�{aJ��mO�&4A�C�&�]H�':m�&0L�7`�S(6�k�uπ��I�������fMBrꂝc@51�.QI,b�{0�9���6�$��^�]��=~0�<zØ�������?4jF���z��ks�0-TG�T
A��_4A��!�ˁ>G頋�7�T�	��5M���P�)L�~�Ԋ0�Z5I����dx�B���A!U�BF	I�cp��t��q����>��ad����
m�������s�/�e��
 `-s�����j_��W�v\|�$���1��n�Eߐ��qc�6���.7�X���"����q��a��I�Uy�'?�g^�$X�v��)��o�-&6�荛�3m��QԤ�n��6ΒА����ɴ:I�$窒�}	#�O��ٮ(�v�C���'�}��r1~�/�>�U�Aޠĸ9�IJU=�z��zǝ��I�k�zs��3?��U�r6��?�M��@`S�c'��,�Y�$N!e��O&;����H�vb��4o�ut8cp�(��9��|$��/�x�eJ �T?4��?;5Ub�b���),D��!�C*������R�[�_{���^��4��:�{"L����#.G̢U�L%MM�+��-������d����u�w�k�r]O�[��߶�� ��ӹ�%��c��S丅C�b�(�O��L��~�q�.����ՊU(�]�����w#7�n�Tk77S.���UG�8��(U����#��8}h�,c��p���kc}��v�o�W8�o�==!g:(B8�sT���i��u��P�ۓ�Mġ5���<`w��^����������_[��Ok�����,; 3�j�SN�r@,��-��)q�����f������eW��OO����$�x�Ck��V�d���w�Nо\�tN.\�$������#%?����υE�[9,�fC��Ñ����,�l�m�4u���U��乌�&�b�`����3��~Y���O��?��4������w�G@ycyE��V��������sM��}�\�`u�)$r �T3yL	��;:P�ܚzL��9��Z��w]���o��ڧ?�6/"5�������~��<�����T�c������.K_������)Ԁ@�j�d�n�@&Ǧ{3#��d��_�xQ��%��[m�U��rDVo��*5�}��ڔ?�˿�`|�ժ�C{z}��mB��-신��sC2�
��͗�v�C�Wm�͔�=�Q�3>a! �O\7h��q�8��i@�Xw{+�i;IT�|��T����lJ�AC�����²���|_����|�#h ���z^�a�]��;�T� �M��n`2��k�i�(��`��m0̄3X�k�"*�pꗭ�	�1�j��ԅ| -M@�77dW����l<�
.����D|�pL%���>6v<�������vJʯ1�|����~�Sɺ\=��Y�
���@�Z(T�bG�U��R��g�� ��^�h"��C� #�0 �}��^4�����;nA6P9}�)5�)��%�":�t�=�a�}׊�j�[�I�~P����g1�x.�.��u��L�'5�5���"���r�>��˯�c?xB�l�J4�,h��c�I��1=��a̪fA�y�E���;~����ѵ*���M��H�,p�N��]���̤�Fi��+����o��p: ��Su��]�����B���R��Z�$�^�Ub�A4�ԿL��=�Ͽ8W����vMJ�z'�����&�d��U����Ӵ��2<���;(��� �!�/�v��	����������,���F:����j*�g$�n��b��u��K��/'	���	�R�Q1��Z�N�-���c�u��G����d���s��%��:�[D��fw�^��10���/,e\��ߤdX�$�ܡ|Ь���NFu� ��QMr�YCYH�đUi��IT��V\��u	�^"�I��KH�M���!W�K���3fx�Ъ�>F����`��>^kB��<5��x<�� q8���j���D��r''�����5]�D�9/�n{�R)���M�bߣr�+��:*���diq�i�ګ�.h��y��%���jD
lۦ�k���ʾɕ�+	�v�I����i����j�^��9*ν!���������~��K�d2�EVd8ѦY)�� �w� �G�'2'NF�����`�C�{v�UYқ$V��� 4mm�3Ͻ ��{�<�������av^��]�$/|범���tH���2��(�i�2Uv,��3z�MS��ʍ�DRׄ�#�~gỏ~W�x����l��ʢ^s�}Lt/�y庬�zj��ި��\�*��x�NA.�NW깪7�7\>H�9��G�Ն%$�M�#}Н9��il^��ռ�{R��I��@�McaE^�|^�}����g��V̍5(�V���%^��8`����	51����6/ǳ�A�|d�ڄ}Lh������Mve���B���A�[ �R� )���wv�OK�zf'���Km�I-�T45ib����@��	y���s��*:4��;%n4"���XMw?��̳G@3��.}LR<�|ygS�b��َ��}�!u�����RC:���MvP���+7�c�v��6�������o��Y��p̪'� X;~�bJ��R�z�n��sݣ~_
~�C}]s�1Z��� ��Tt/�&�g_�I:��9���ψjcY�*���u��`�� ���D�;��2����.�CUq����H�D�;5YXt�B�M���I�������|�b]����T=������L���&���9�zc�&z&��.�Glm^���5=[�r�@�b��Ԡ���r�V�2��]}����X'��h`_�r�t}{[���y:�L��'z,3*}�����*�c �f��s����b��9LOQ���wHC�8�؊Th;c��6���z�(o(Y�:cEV�p:.=���2�X���? l2��x�Ц��yHX���`�x�É�2_�?�d�f����O߄�������mBG��E`��o��F�lJ�?x��m�ʇ��^�p+y�����j�0챵��#7����V��6f�'�*����%��~:6�[^��ƼĎ}~�p �;
>b[��(72^C`D� ���B�f�Zh?$l-�,7s��;��zV#8���H5�����Mҡ���Z� ��P���,�����,�u��Tp13f6�|lY�E���Ln�Z,E�G��]>6rfԳ��u�x�\���˞z#�a��}���F��-�>�}ii��k^߯:?��@�ȵ�-�淾*o\Y���N*ѕ׃��0�v��÷�ۼo�����߽���A7}楈�q��6�{����\	c�B��g�1h�!�Is�x"'�����d�"5^0�}�@���85� O�\[5r�� $�:� �S</K��ԉ����/���=s�Ѐ��<��:Þ�.4����ۖ4*��Rm�X�'h��@�/���P��g����� !��,5��lrZ�Z���н������˜ ��]���r�ouq^v�ٺ֒�:�(�9
L2�p�����w	}'ª[$�Ӆ+  ���3Lq>��;�Y]!Kg{C�X;+G��h��>~����'�w�M��r�l("�;8�vu:w�H ������Z�̮ gM7��@B`D�l#'e����n�Lab&�f�N�� ;�Ѱ�`1+BkGF[�@etX�v��V$W+?��ι������.JU��7>�9�#cV� �0�H�<�Ŀr0�k��9!�:՚�s�I6����N��m2&�P�q��_��ݝ1H�彑"
Y���A�)`&���OL=d�j׮]�/�V�zFl�$$�&��ㅠ򌝎�xX�D �{�?�}�:hUWY�U�?E'� {0�\+�;F�'3�Rǧ�u#��倡�>%�ҀC��Ae���r�z�aɺ-LVLX�heR���v�͙�U�b��RDr�ZteK�Ɇ��^;'/�;'ϟ�,k����e	4x쏐vV�^V[�j���#���d��� �����x��� t�=�ng �.����U��\�ؑW�</�;}ixxAmD�o�:�K�W���&Vt�qJ���b�N�uGEV��L*�DV��ĵ���d>���}P>1�<��!����fm^_���׳�Χ�[� [�C����	�هĈ�6��o0����f�Y�+;�= v��H��p��y�������L%����t�"4m��/_�6����_�t��kp�'J�ƪ�P
�r�&��^N�����W���k��'>"���f����r�@؝�*�X�-������j_%�3ガ
8�l2�f�6��C짭Y�33L�؂u��U��V� �[�n8g��C�ޘ8G��sVh���m��U�3����44���8����9t�;єh�TV�8�$��=kZT#�Ɓ@�]0��I�'f�h3L�s�:�nMM̈́~�����.CϻUNXK5�|�ZgƉ���Oɥk���>�l��瞓�?���_�&�ƂTUg_�������d�}�~�W�9�5���_���ԃSx�lB�q�y��K�OLÁ��:�TS�T��;�^�\N8]^�̑2g�K�����pA�JSϪ�E8g#7��ϕ�-�ؑ<?��
x�t��_<+���K{s]s|�����'/�}��C� _�ܑ=u2~ڃ�A�2jk�֥MmSE�\��C����֬�ՍO����)B|xaYנ+#WW���S>��{�J�S����s�ț�.��g�T="&��4��4�YVg��HVR�sw����'���s�ο�oG�������4J�Q�(^�@(�[N�!w�~J���r��5���R�'�lE����58�j�;617'��ϭ��5�I�=!��������}A +�(IⰋo�L0�@���/�<"9s�t\�v$U����4Գ�� i�,���l�D�G��[۔v��%y�g���KW����~�)�yB��aK~�@�z�!�+�
$��8r�>ܴ�58��U�$�4� �%�ȉ�kU��F�Ǥ-d��U�p4ƫ�K��%��	�f��U�}�?Ȱj@��ǹ�p!�\m�P��b���`җ\�8��tt�6'��w� ���5�[QrP^ \��l.�z���.[��p
Å��Q���S�`�п҅j.U���(��%� �����p��n(&$<�`��3ih
c^�øx�m�%Olf(}�/�Y���iy��i ��5,k�5�ę�,����&j`������)��n9�Tߡ{��KK��,nV�h���K?��A�J%��n".�%���S���o��i�y�#��UI��uE� ���v:�[R��]j	J��pWHo�a&�P�Gjr������mL�2P`�Tc�u:	�!;�T��h=��M��J�#��O̰��b�-��=]p!����ӑ�E),e�Q�F��V6�')~~"[�.PW�	H�K��Td�\�[�I9$����&T��$5����Jd�S��q�;8`)!+��IfأHxH0t�ڍ#�k�__Z����'���[��n��r$���~���	����A���"B�<��)X{s���:�;{DS�S,��d2�3�G�PF.W����Q�eL���31��M�#�M�h�&�Ӡ
���qYQr1�s���#��D\賽��oql�l� �L�nJ#T�\p�/r�
L�⏟������rx�2l y٧��3�J�$��iL�[�@�3$�uez�wS)'��ep�FF����@�.a@]ҽ�D '�G*�z�{�����$����D�ly�V=P��(��㝴Vf��y��E����'��%���>Y�;m�n���l��_��G����D���C6.����RA�hЖ��u)�9ih ]Ǭ6��1���xе<��ϥ���g����rm���k��6ݫJU�R�� �x�45ȵ�`l�١+A��~O��j�$G�����n�uN:� �!��Kس��5�d%F��'�u�|�C�#��C���g�����ŷ��e��M*��ElT��c�	�Ss��c?�U�BRЄ��Ҙ<I#i4���!T�W��j�u����ꊼ��w���,�ϳ��s��{��ʫ+s��TΞ=+z��{�]i���y���*r��iD{u~���U�9��;W5YW[�6�hsA��ߑq{[�ߓ[N����㲀����{ߕ�������ȥ3�58lIY���BM�t�G���	�HФ}�re*B���$4�a8@L�/�]qH��'e�r�j��� 61��`#3��D.��O�T�1N���>`�k�o� �m��jZ!]��,'���礫g������R[�Z]��l���@6��(O?������{����λ�һ����S'����F=R����,2��abRzV97~C<�j�J��8�1�SW!��NY�dҊʮ�_G�
-s�[��\Az&��m��ɃDϥ��.��C=}���Y�Cek�$Np$���\߶�.���F��M�@���Yq`��$f�׵�vj`Th�2j���Oa�����!l�h���7����'O�u�����Y��_*�]�u���{ T@�(�������|B�?�P����8�C�(e��������!���4���J��u�!i���El�3��puIᤧk: �?��qܧݘ��QI�[	�-I��n�O���D(��r���~�rh�"_�ޏIv��
/D`r�w&�Q�ȵ1��n��$����:�����FC�����K�V�Ej �֮�YW߬$�8�kV�:T��s�����Ij�X��g4J��U��
9�i�y⸓@�cD/$C�����5����y�М_�SRC���,i�X�b#g���'u�7���X.��ɛ��ə�oIk�-M��#`Ot��9�l6���A�	�X8(ui�'��Ar�rL�i#���>&l1V�vk[���g<��Ɛ��M�,1ohp�!�j�Y�g�R��.ϼ�|��=w�����p��wc⦶K�2�V��"��L0	��<Zh'c�|�̀)gh%��<?�M��ڴ��=L��Ij���������&�����@]uj�x�rb��e%N��J��clT1��=9�p�]��Y�ĽE�&�֔�J�'�i��eY����2Ht�(���\����{
�����n��I=5�.�-��8b�\x_��?��y仔u���	9}���e(�,��X����Wb�:'����Q�����./�Ƕ���7���*��@��PD�*\S�礽��$굥:j���>iKC���}�~��c5@h�4�^�*��p��J��s,�))���I��(�@���04Q�n�X5'癇=�u,���/�>�������{�v�ˢ:�yu���:��A���@���^�s/<-W�(sPlI����e�����f�]Mfd�9D�F%�Dw�df�-�� ���`���@��T�D^U�,4�Z��dqi����
y5�[�!���1�k����Z4�>�X��fW_�kW�3eE���u@a��]H=�Y�IFk}%�r�D��P� i�ɥE����ۓK�^S��#��8.��؇�8��^,��,w�vJ�j2Pw��i)�=Mu4�@��;=��v�i ؕ��1:�BdCc�dŰ�>����Qm8� �g�����wv?N�*��%|؟��d� �$b$t�2�g9�g<rvK�_�50�	R����Cpb�%U��u�ww�5�R,W�o�!�\�,��8!����u�I�i�|��Qw�k"�iQv��X�b��F��aDDtk2���`�A�<]W��r3z}'���5��s���$�.T6�)C�lR��dc���՟��w�]��`��Ѭ��{���%��r�{�v��`n��,�1�<)��R��0���U���5Ҡpl+L/SO~�������ь��s�����k�}�á�Ę8M��T�ك�((��s�49xAֶ[rU��!�!u�P5�/tp$g�4ɦ��D��{��,�ט@C���>����]_��8���g�*��}��I���Уj#�[�i���w�����Y�c9�=��9YQV�5&��p�ve��J����˱���:v���R�(�&�����r74�x���<�\��nG�w~U�t����p40�SZ,�y�P�$aj�7��Z�G��>�b���h�鶑�^7,�n�+�ww��jMn9|����[�&��eZ��b``�j��p`��a˚!�q�.y���o�ɏ~���ziCv��:o�Y�[�V�|j��~B��CQ�����~Ǹ��-XC;� PR�[H�Љn��8!�&�[���=N�;6�JR� �MP������|����֮|䁼�6���4�J7M☸R��g��+�\<�Lr+���4t��M
1��3���3,� ˪����Ye.e���@X�IxBd��xl����zv��(C�y��(;��J.�����a��M�u��\��m��ShBG��vs�}f��)�佼���#�A��%��hA�%2�S(�t��He�Űb�<� �����C��_��<��T�9X�5�ȉ�rm���i�6v�N=IG�fi�m�W�s�k��y�����B����i�r�Q�lүK���n�Af�u��XAA���$�Dr�J����C׬�#G������w���r��	ihƝ5S�kB��k��Φt�|�yἜ;}^�}(ǎ,�����:�ڋ�rA���M�j⪊u �um����)�;��Y�ֵ����Tӌ8�[N���~���p���A��\�p������C؀g�Z�4�)�%�� #c-p�>pn@UGTe0,�=ؑC+�2?���-�L'���:w欬���#9"�EYZX #AC�^N��xoO��u�S��l�id�w��F�yh�[��$����?`��gwgMz���m��%N>�ll�֠K���'��{�'��yJv0���L0%���)kb��C�z�({�5���&�W���f0OB�Xz�K�9:�b��E�Jk�9I� 7���y���Y��fA��.��d�\�wCcR#�.ML߸���I���,V�%��P׿�{�Hɺ��"�ku^�`�t�V���قVP(�ݝm�|�u��^�a�Hu��>�D��%}��>�]Y�U��w�'��*�9�;��g�{P��L�al��٬Z�������%�}z�C���1���'�%���<���$���@dF�H�&�1_�$����@�>���H���=fP�!�<� 5(f�ׄDg
BǬa*�bN��ϖt���9PCm��ͩ���-�$�R���:b�І�pϤ�,Sa-4%�|���5��H��a�N������\�,��I�=���"*թ����,&�3����Ne�1��`E�w���e=���X�������s�o�^� ή&�C�W�������&����X����w����~�ye}S݊�%�H2��8���P�Rܓz9�{O���q�]lj��e����\A��@Z�Hŀ4h|�M�>~���[���Ͽ�k�\T�]ԯ���Z�^�':q��b����Ś����tms�o�#�(r��n�#+���{n;�/ܢc)W0�`�Z�u�W4��q2_�.��y�a����)������޸ k �"8ҍ�cP*4��ć��>�_�׎�7�hE#�~�c�B�����je���"�s�(O.��A,_��w�ų�4���&�pu�p����i�	&�QE��!]���tV^~��wם���ڡ���t�ϔ!ק�S���Ѧa��x[/o����r��4/2wJ(�L0��Ye���V�7c'�z�Il� L&�x����,s���Ft>4H�L(5*����s `rsCKY�%D�q��)gW	4)��H�%qj!���:]iq�vb7�ű�Z�?���i�z� c@�T�����%��Ꝙ�4�6s,}�v��e	�
v{c_��$�Bm^���7�]��r�2[	a�DC6	F����S�׬�������F�A�����tn�W}���>��CWID�XH ��� !a�+��H�r�;n�O?��T�0�9:��M���cG�	�A�1'��D�Sg���"W.^��9ҁh�8Le�5�X�O�V# ��o(���W4��JU�Z��޵+�1�ʝ��*�;*��s�ɏ� ����eA8�c{{��ۜ3iK��v4 @PV��������ej-׫s2@;+��A�<�6�JT��A�|a��ƽfS�\�����%=�e��x̩[o˜r�a�bbr'ġ9���I�Ԑ��@Z=��_�������c�w��Txk�G9z�,��_� Ľ��G-�C���=�*{;��8;r�[�z���EJ͡�k�e��mC�8Kz �)L"i���}���34��L12L�$5�)�H3{���V����V�,��,3���۸H�щ�����5t[����%ґ������ۡ{Y���Z��� ԼA��|p��@]=�mЍA�q��@@C���M�����$n�ޒ�'���:��~�!���,TL��CP��ʦZ*N?;	�'L�Ǳ��t-�@�M�����l[{�k]������6_-2�C`������&b�ed�9T�@�8I���둳V�&Z�G���ߔY&��!X��Xb���"�C��0�Q&np��?ӌ.����]�)�?�cj=G�ْx��D(,�1�'|F��ʝ�$9�(t��h��#I�8�%��c	��/�K^�pI~��'Y=.��HP�*:����߃���f1홑�ZΡ�J+�y����ǟ�q�*��C��%�k����y��{%Gn̷����lKV�W�=����՞�5��{�C����ڃ((i�X ��f�����X>��w�{o9)y��y���y1쉘A?� ä��&�t[jÁ�nK��{��4�}����^�����]ʳp
1� ��L�F2P��(gq��M���l���U58����?p�4��D$ �U���cG$���V ���uẝ�t��Bk�j��7?�a�瞻�O��\��Sn �
 �<>����;��⹋�ج�a�qZi�J��[j��n�@��P�x1��(��/��^�X?��:W�t�.�׷��gȉ�d��jY��0O44��u���j���kge�՗���8u�:��(Ui<��b�@W�863|�\���
�EIM��x�"�����C��pd�o���3�5a�"kxrs'Y��@�пī�H&Ue�;̴)�n&�~ׂK���eX�BбU�o&	�+_\:j���괵2�p=u��>w���G�mk�p��d�k=	A�q�^CV1��c�&��C�M��Z�����V5��~m]旗dS3�+�a>�����^S�:b�p8J���q�K9���@�G��p�o0�f%�@�9F��W�*�6m��!�ך�h�ܣ_��~хD`�/���=�������8р"��y{�.I��J��=�=rϬ���74�FP E�3:i�#�����3?A�:��4����3���
�Zݵt-��{Ff싻���YU�0�7
U����={�̮]�1�g_��|��_���Ľ��2�����Y�Z�q<"(��g�9=&��Uȓ�7<��`0�&��ΒzΗ�~���#cY�|]�pSx��֨�?)HI���JK6Ա��Λ��;��z�m�׮\�����*� T���SԿ!3�{AJ���=Fw0/a�767��^֥^�V]�{e����o~�5�����ֽ9�����p}ӓ?�N7ڂ�,5�ʥMu��r��]���*5j�[�N�a�<��K�̶��<�1����>::��M��t� ���'���eҝ��gR5AY��5��M��_G"I��t)����$W�����]��;�����ʆ���s�,ҪX���
�P��XC����7����2�t��JeټpI�v�y��FŌ���i�����]�rc�6i����Q[�|�fq2���窀�P|kS���%�f�O4��z��`]�������<���T����&H�0�:� @i6=#�!2�^��aSA��vp|(�nGJ��4��]n5$h�9E��.xm%l�hKD�����<���uy��嚂-p���{�P's:��rh��v �'��Q`c�]˞'Q�Q��f��|��lf�x�K��y����;�l!�X�d�G�����p�����u!�cZ�m8ZaR���iC��'އ�'@��#[��p����(=���Y��E�!	����	V��-]u�"SŢ R
Jt`����3�P� �p#��j���(��D��$ۊi��"��D��j�#L(x8%_�Mj]��=�O()b� �������?�so4�^�rv�~ڞ4�6d �'�$$-�^����|4����7ߗ��/��˗y�Ph���>'wչ����Ȕer����sq6���K�_|�Yyn�%K��rtx�!Vۂt����u�JQH >;�*�ۓ�n�b�����?���R�eO�~禔�ejm"�7F�S� �XH��ĝ�������cYj�PW�Qo��5��!S8���^���%�Dc�XD�X���&HC$�� �V�3��V ��B��4��CDs�7���%���#����{��	w�eY�G����Z�].N����Ca���ֆ�P��H�Q!�d0>�r���@�]�"�HUlL�a����myW�%t�bW�|�H�8XP�5-��+X�D_��ݣ#���KEϽ{|,�z]�U� _�XU�7*���]��B;���*�����ĝ!8W��8i�`����nAH�-TL[�D�8N#H�K7����Ը7��s��O�=�U)[
 �1O;��ÝYu��n����N�sr ��{�s�(aRd��1�y��� �:h(�^DN��oօ]b��U��L!���a����/�e�ZC����O��;�~Dg�C���6qSOA�N�R��x')qK�#ZKc���IQʯZ�l�u�_K����Oe���jkf�4��7�� eA�{MǬ�0��	�d��_����w��U�>��+������Xڒ9r��ԇ�?<���7�b�`//���ɩ��T�����כ_��r�#UO	���DOe������W<���e�\_�K[�,v� w�6e�Ϊ�ں��	h�����щ�x?yȴs}yC�OU�V�䓝#9=9�K��{��;���PNN;�`V8�id,���Ez8	)����4rM7&�/�fR�.3:N"�'N���34X�6;;뱈`	�r�~��V�����ҫ����R�桶�M	(Q'�/��I\�ɣ�{�Iɚ��U\5�W��ū��A�y�XaJ"2u�WV�r������a�@JZ����u,`�=Y�ԑ�uvzȈc����[A�d^hY��9x���s�H�'a<�b� �(0SUu0Q�<V��+��h�� ���D����I�U�D�vTDU���JN��Xb��J<꾐W�_�ړ՛۪�HA��б��Yұ�P�ⶼu�����{૲��Eɥ:����Ot{]�%Ω"���_��Sq|Ϫ�1��20P���jK�u]c���8����C�=�13��QJ����D��*�{�e��z�7�x�M)J��͎�9���T��M�D�k�<��G�85*�X|�ŵ��(�1�멩���S�ݲ��h��s�׵1�����D^�=y�"e��#�Kc��u��EL;Hf_6�T�Ӹ���VxcOd1���6��E�!���x���پrϋؖׯ��v*��;2P�ū�ض�s2�2���ya�1���L�|��k�:�^Om�8���K�Wk^�ZS�i��#�>�j����px���F������|��<�ʫ�~��,�z��e��3j�#��QE�v����^/~)�n4����gނ<���ވ"�%5VϮ5�w������X�/X��\��TW��Ϸ+���]��g�R�]�8����t����o~�2pwV�E]�we}���7�.����/��p[59�ɿ��?c[��~�r�^���	�
u�˅ա>$��])�Q�XG��G{�������lCVt�a}�[r�ѡ,o\��b��sG�^���.���6yj���4�0I�[j`���믾"_��WusYQp|*m���,�N�_�h8#��[��u��Y�I�`����F:�%zf_dn(`�C��%i
wz�Z���ؕ*F.�k&]%y�M ��,1KZ�]'�)�'E�sab�#F<w-A&5j���ACH���?��uļ���U*���yܤ&�;`�*p�r�P�5Y�*�YZ�$����Xn޹#w�=���5�9�"��QT�,�Qq��D?I���N�X}�.|V<O����xJ:���k�����H��w�	3f�ʐ8�E2Uc#����R� �?{]��vA�>`ǈ�Ֆ���.�!;����W�\C_j��t���$ѣ�h��H_��;ݓ�>��T��_.��JWR���)�b�z��}V=�݆��y mF}QN!�S(��XZgk�w޿E����>l�}E�g�N=5�����e�=ط��>0�����(�!5<�熍��}�Թ�	�:ꍪLP��w̴�G{�(�Սu������K��\�Q�D���1GT(�б�)b��͋k�?ұ8:�k�Xp�=!��P����x�#�-��:�5�v��esu�ڂ�Pn\�&/|�U���Er2���E���A�Z���(��:r�Fz�EF$B������9�#+�4-�ɵk�3�2�{%T�E_';/ӵ��I���Kh�Z���z���]aC��6�fC��6�k��\�K��n��y��GñΧ@�z?��ٰ	
:�T�h�ɽ�:��#�@Pd�Y��7czr�7�9�MB��9�ݿ�����o�ƽ"_A�o��o0c�E}�љ��oٚ��T,V�ik�U�z	����lnm�����md��µ)����9'1�K=��mD��7�|��E�cO�O��D$�从_9�i%3�`�H��y�ah�v��)}�6D�.%�g�/`_k�9+TAAN@�~�{\�3���c���jW�a��5(���row_��w�/��4Nt��x�?���֔�>�����
[(��>W��ަ�H�\g5��x�w������>��2��,���Qsq����PR��^���۷e2<V[ٖJ�N1�rP� ���Ǟ��Օ�|���ʕfAj�:���륲4Z�P��Z@��ڌ̪��N�J��+�.�����m�}��we����y�YrpQ��e t�����t=�wp�)G���;�X'&4���jT~��/ɖ��A�H��"T�������R���R�+��Vc�+���*,�M C~��?��{w��ɾ9le5D�RN�ܑ�����_��O_��j����������w��I4��=��'RӉV������we}u���2o���o����z�h�ņ�2cZ���E��\G�uS�gJ�L5<�k r���<��w���n�%ί��\[k��ș���qF�x�{��O½�);	�(S����C�n��Ed ��Y2��4���u'�{J��F)P�1�9�X?����\��|����E-'���w3x����8�/�x�Q���B䀫�M�'�:��L�F�=@d�+�)�9.n�t�-�z��Jw�B^������wt~�G� L[�*������b��4�h<�)HM����|��J�ؕ�ENW���[ ���4�|�Eq��Q�t*V�)Gzn#����JQ��P�ѮT"H�Ĳڬ��7�����P����PE�.-t��1����#i�׾�n�
2Tח�%ZKV�2�ŌĠ��k�L�Z����c9����{�pm��JS��wI�����f�|2���M �c����}���v�^��x��$@���2t�ӛ����ǀ|i��w�������8��ov	9�,�^�Nu !�bm�p�6��W�4��W����t���C*	������ui�k2S���0ꁴ���K7��I_�����J��p:T0���YoS�stH.z#�RQg�կ|E7��EyF�EE$����ܽ{�xT�sVl-�>G�<�G��g�3�H, b~ZlńQ�1�ZR�k������lC�y�8��Į�6$4
PP;<Fj]�#��u� j����� �O �޷�,�)��]@Jk���#��A�]Ag8���33���ڹac��2�����(v�U9�PAL���Yo�H�s��7ss{_O����ޕ�����;�\^�~�X1i��$`�u̲([�v�y�<mL���~ao]ز�葫7�#�?�Eʪ�']��Oa��w�/Ra����O�(d����Y,��J�!p1�w�A�GRh��P9�9I=�'س!�C�/��Q���Q�Ae�4�uǥlqvD�rlW�l0G��)-�ɾ:������{��;�R�4���݆�j}Y�?d!P��d�� �~4xwv7�D��|u�QU���:�ݬ+-�|�=��y��jŋ���Ə���V������:�����9-� p���\V���:K
FWt�^X[��E���0b��f
VLmSEߴ��\��^ek]9��Cپ��T��,�(?~�]u6Glc��8ޘ�"�l@�<ltT����}Б������ɳ�ٌ:��2S���ٔ�7�����ɛD���(��Jf�ɴi����r��������{r���� ��xO��e�ҵKr��Ƀ*U�e��B(_nH��  �`���sWn�ߓ���U��}�2���}9QO]oDw��P��F��\�����j�/\hGd��@��t���u��N�nQ��������=y��m�ݯ~Q~�K/�d��鳜GC��A]��y#���i�f!����bJ��� ��{>՝�-�w�Hϙ�ӡ��h��1����7��A�ς~C��	�:Mlu���)�Q6�;�^Zv
&p-CX��<���a�R��Q9��m$鸖��鑼������ӎD� ��2S�nF'�q*�n"!D���D{�)*��:!Sg�t[�����<y �Xg�.�b�3��@��	�}���Zό��v��7�Fb՜q�4'`0�t9X�D/�q����O��O�؎;�j�� �D��48N�e��+�5�;x(ӳ#iVLzdcc��A��z6��非|�s��f�)Qo"�oݓ���Ѱ�b��e�,��y�}��8�:H{�� ��qƲ����gё_�浫�Q ���!�q�+"�s��i��QS�UD;ET���p�`�CpG���w�	~�y�F Tk�5xN�*F�zUߨ��ua��c��c����bh��S�0Ùk*^U��!*a��8 S�u���+8�� ��Y�!<���UF����@�6۴��:���7,(�]ؔig��ɑ�j��M����3�-�duu].��\ZF�r*8^�7#Gz��h�D7�.+"1���%�~U�eg_�.\T�Ґ7�|[�����js�r@�#�UNg�sʴO�Q$rD�J��,97_]{�8q^��J�~1j�OXM�.���*�#���ؤ[�	����O�\�{��Dܾ")yDGuN�[@��"I�+�#{*��YO]F��6CZ[Vw���F�\J��+�L�U��D���'�ݝG�}y��E���肔��\[H���.�  }��\k;�P�Q)A�����"�7���E�X�)I+�<�F�$t�c8��T>Ƥ��|�8�2
����LD6�ȖY��Y�AH�x��8H}���tKc�{�22��v�M��=u�F:'�KMf��~��g(+���`��06�D�=@p�7��޽)o���쪽��dU�S@M�`���9Bτ��Z:n����Z,�rA�a `W��R��������;W�I_m��Eݳǡ������4��^.����G����o4)(���:��Bʏy�A!_�,���M��(Ȋ���V�_�#Q�(<q�C9{O�Q��Wl����z
0^���4�;j\zNs  �AIDATGE�cU�W��&��?R�L��-����������� &8���)y������uw�������vM6���/�{�$��z��[�-L!1�k�ȳ;�j���qI>D0!��zh/����	7kuw�6R{�I�������/��Q�ǂ*���}����z�
2u��xH2�cW����	sb~X�(5�I�眗��pS�L��/0.⮂�����;;��qaU�6W%���J�����n*��乹A�*d��1���bya�م�A.�J��y�I!����'邀)\�L���5��_��AZMm})����h�VV����u��^�n����9g��Q� �ɤc�:�Ď��k�K��牥�CkRI�{�V4�y���i7���������M��?��Tc}iI�kW(�nYv�So�Q�)�m��^1K��E�=�u�p��,k���*�</��W^Y� �4�iEx�[<�it\D�U��������О�Zjʕ�˲��FC�(��k��ցz������Y琲O�F�\�{ߦ�S�Y�~��g����m8e)N�
8�\^1º��b��9<R��ho���H���U;�R�"��tT��>D�@�9�ݖ��쮩-Z]i���\�Z%_�hG��Z��FN���>�l��n5�K�%9>:%]#i���"e�n?톂��2ub�ձ�B���I��48Ne]�H�A�`@���뾞�P�"�,��t�o
��nz�mS&H7�cTt�:ᙌ�=n�����}�&������견��m�X�k�ɑ���L�i�ƀ9� Y(<#�j8%?>�Z]��+�+5�6� )��գ��R���)S�Xp�����,�~���'Z�����N�O���� ���<P��FK��1����tC�<��Q�pf6���XN8G=F�����S�4j��k׺��if�Ow �K8M
�+
*Ů�y��̳�Fv��k������rEA��_�����3WYu�"���uiOӨ8F��p<3�2��|��$��o��Q$ݵ=K#[�`@R��B�\�'��V��'�R�FJ�!�)�7�p���G��Z��r]P8a!!���\��"#�x� �oAp{f�#���������8o�l��(��K�T�<7��Q�||ܕ?��woߕS]7���C�u��H�z�e��Ա��*sw}��P����SҨxf���W�,M��*��L:�Fт,��wUӶO�q@e�؞:�aƁ�V*�Xg K�7d�ҏ>>(�t_�����,W���������v+y�ڞ���x����^���4��|�v-7�겵�Vܤ�:(3��.�t3$���Ōih[��|Q=����t�誁YׇwE�c���1�Ip�Ԫ �t��Ȼ������Y�B��V}�\{e}K^����c��b)LDzBg���"J�l����2� z��C*f����J/�̭��A��>����Β�n��r���]��!a��@�E7�\�ț�o������Ez��E�?��ɺz��j]7"5N�e�(H�dA4���.�s�`�� �EN񉼏���Xa%\hdL1x����aa>/?��q���}R�0dE8���b7t<)6��ª8�C\�(R$ ��ER0��q�w�)��'/��̌�����i�~��^τΘ��+T	:^�w�Y%��{�O���Sn>:�����n�mT����ES�̀i�%H8(qL���@�2��w'N"���}�D�=��Ĺ���	�#x�I�$3�� ����N:OS�祟[�}l�KY&�(X�Fj0b*��cC�^ǰ3��`(9�*EThШ��?�~
���CK�����)+�+�R[]��u�v}��f��Ҁ辄��w����}��6��� �����}:c�
�8����@p�O}�uݬ9ct�y�-���ԵV�N)/͕�pV �'g
B�N�V�ň ��|��w�~���)����)�`�M�F���A!	�'p��v�<FN����#�Q�7�Jby�%����n���*	H�kvj�� ��"�� ���㱱���'�n��c�+��~.G��p<J�����7
��@� U���3
3���b�.:����؂�Q�ٕĥ�9N��w�o4��E4�$R�-e�?a Ϥg(efڼ8��Uj꾃t!ӷS����l`��9n���P�|n��A^�Dduj�L�)RiP'�H����;�eL�kF�9k|�ɔ�\{�b�,���z�?�q끼}��\�|I*A,+���o}CZ�25,g:g. ����{s�MF��'�X�	p4�u+��N��Q���E�����m�Z����)��B��`H�g(A3��2�hV�YUw�x�iw���lD�0�y�Ո�B����ZSt4`��G@E�X��QO�}Qm5Z_޼'��<���C�~�'SWG�:T��=��!�����l|����KI)9����}?�0z�f�"�Y[�(Đ�1s$��N�TW5�SQ�W%�����#��:�쁎m�m�g,��ҍ��b��t��Sݘ��O�NC����i�,k- �S�����?@ƥ�/��-yF�7�[[c~j�^8�#�d��!�UE��K>�ݕ���C-ʕ7��_A)�Eт�]��aR n1�$\�X�2ף;��z�����A$��K^+U��ȍ��7��Ⱥ� �X)��,���y{���1i@�F�2ѱ��������"�|>�T.������t8S\�X*@i �TnPhv�JKz�������+[����{���V��y��З�=o��j�O���Y�s)�{���@��%�Q<��-�A��%������62�X߁rUPY��"� ݘ�'�����ZIWT>W��͈�Y��l���v3�4�Ѽkdj�(&L�XQV�Wei}����$_n�����-���]���^�n��ǡY_F͜�EA�^��$�e���֛ڋ�|�%�خ�3��ӊ�d|]ڧq
��g�.>f��"�8��3d���)�=��#
t�"Lg
ؒ�ĉ�gKĦ�8G]L�MUA�T������}F�PHq�P���z�����2�q�Ξ����
\�HzNR�P�(�����͝$T�^Ӎ���l���Lu]`ހ>�u���D.^�(�/mq�S�{r w�=K٫��'�i���T��Dm
����$�G�a�� R�,꿧��ʁEѧ�T���_]�<8Z�M��v�L٣�Ѩ��ޮ�G�1�[�T�Sc<P�~��$�| ��GBC��+�Xg
�����3YZ^�K6��Ɔ���`���7�GqD�q���At�/i�	6X|���@
JA@C�i9�m���b��Yz m���E%	+f�3�6&ݴB�6�Ȕ^lE�}�%(&l��W�mC��+ ���v���i�ƕ!�����D��E�Hw�,� ��׽$ʌfE��Q�bS�k�WjX�v��<~�x~���(-^��ň��3�Z����~���î����֭�������%i�ܾ|�9n�ӣA�4H˅��JJ��.@� �oE��P���t:��o�r��wƔ2rjxt&�򼉖m���匽��(Tf��^ręsf�[x20)��p�Q���uQ������`D�PE�cgt_����w��<�y9�{<>0RX�4���,�Y����т��Zt��ya��1C<���i5�m'6�?��|_�-�ERĂ�z�� ��M-�2m�tP�2g���gY���UyB�ky�W(�2�:9�	��j��NĲ����`2Q��F�}�{͞I�vb�X�P��j�Cs����*�G�V����\��/�Y���T�w�,��՘4���B�Q��^x^͚g�-s���9���t`� �7k2>ؗ���ԋ{����������w� �FV,I&�R��[�b	h�#e3��8!���ލ�� ��d�%�'<��
3�����>�䛆����������|��.�������X���������]y�����"���\�ܔg�^�-H�\�$2�M�T��G=�)�O����$��u6�|�-�=����"5��A�ʫZ�%w[�ݠ��w���&�=�:d7�ڙ�+�4���fLmY�ؾ)x]�tOD�ً�� �n��ހ�*����"=��(�.fG7�׿��e'�;�w�[����7����Ga�H�,9�Q���*�0i�s`e.9�|G"q��Rb"�I%r�KS��%<hv���8�ќ(���$ �ˤ��Y�{���$��%�X���n�T��r3�ABڣH�+ �V�a+Y�,v�&<9>�g�_�/|�%nhu�F%Ov�N?y�Cy_7�:4�nݞZ��pV�|V�A+�j������]/psΤ��L��@=�B����ޑ��#�>�)�.��K/=C`{xp�9}����k��n`O=�[���. �r�!HD��ʕ9��I/u `r�i����v�^K:����̵�츀���'G
�N��������:��kc����,��~p�:e=�+K-�څ����M�vj��O��N�Hm�z�(f�����֭��l��햂�
��_v�R{s��\D�0��)8����$���QGn�����'U�����M�*P@`��WC�􌽎m�9?��X�u��q$�Fj�zN���d��?���hd]B��Mק�:� 
�t2�Hp�v�?����]��G'2�9saiY�Y@�l��^�?9%
T�r�Ei���z>�U�uc�G�p4�,P�=/�[�Y����#0�(�Qa<����h^�,������?�N��?cC�F� ��xF��ҋrqu���0��>���w}ƿ���G{]����P<�w��Q͊O����FIPtf�C�;�cO�vN�"�cd��nR�� ���,vB[L�?#d`{�+�����3y6���hu�Tl�x�����޼��q�ǧ�F����e��ޕ7�~Ou��YI�ʾ��	{��39���F����}FO�%�i����L7 �<�c�ņT%���^&
pN�a �k?��^�Nt��!��������Ql�'ߋ+�-U\(���uǚ�ە�_Dp��W�0���	\UǴ�A�Şl��\�u���ܴ�c^�m���e	=�r%�N��y�g�8`P|�pX'��<R.Y �f�� �2+
 � "$T��E�n�����5�I�����Z[���jH�j|�e�z&+�CUmq��qF���dF-�	=�{���L�g��d��F	ùn��q΋xj�?->�����f
�b��B!w*���9�rs]n��M���	�=?��u��s��o}�+��l!�[+���}�1=�[ā��7Y���
�6C'��������F��Y`�CW��%:Wֳ�s�a��c�g�	��,u�wΜ�k��܁�ȇʛ�5�Q��CT��ρ����H���Ρ��_���~�C�NW�'�g��V�~�:	������Y��6w���;	u����J��<`��7�.NZ�%K���#q���,P4nh,���8~ir��)j8*�L��AxU����pm�ޏ"�j���*���Þz�G�z�`d�`o_��ug��_�|Y���}x�FΎΎ�gc+ԚLL2cD6��
���1�S�x���N�r�V���+�R.b��,F���9�Nt����-�C�s7� ~��-���1W����dgg��ې�$WR{��	7j
�3��P6W�
D/ʋ�?G>��������.�A^�rQ�g��� ��� D�H;��M�iW�\���e��X�hN&5� �3��� ��0p�nc-M��p(�P��9�9��Fp� �z�y?`�?������'FG �#��?�S5���
M���̑��(��Y9�5���3�:Qk4Jw2�;�Ǽ�qצ��A� ���Sp̆D��s:��.LX`�g���r��-�LFN��g����
�8Ƕ�u�l�y7^2'ܝe�Y�`;6z�s彺���X�i��i��4_�J̾�i9��L��~����[��f���x"�|��0��y�/I����iGӐ�2:A� �#5A�+���`�^pΟ�Z2m�<�a�Hl��6'h�J9���^��uѬ7\w6�"��lf�v���HQ�L���2^��ֺ,�~o�eJ�ܫ�PQ;��}�*���&�ư�5���C#�r��?3��A�ob��Yd�=�%��=sD�siZ�U������*
�X�8�Z��iu����-�S�9pp����B���:G��}��%y���^�Y�� P��i����se[E�Ib8�������~2�$Sh?z�z;��=GUdg�%_ΰ�GR���="_(�1������D�nO����U�&�׷��g0^�$�����#����C�K��t�t;�-�������,�@^��\���^���V�IW�!�j�Z�{t@���Z-n؉�h��8��|�$��髞�,r0)X�D(���?	�¤8���/2�ʹ�D�#��º*u�ȳ|����sW��o�A�T�����M�Z_&�r"�-��B[9�"��>�=\�ӸD�c�U�a�vr��^�w�2������x��JQHE�ߨ��������������<�c�ڃ�B�e����<���_� ;���Zca�����W������,�����~Sq�2{v��Ⱥ� �"�p�%��<���a���9�C'�lɞ�9�|&�����yNS�={�<���a�����!f�r6kTS?3�q3}B���
D�0�x �k�/����`ZE��H�֖^xN>�����DlPH7�t.#��h�37��ƛoJ��1�_�g�DB;t�`@{�j�ȁD�Qs���ɣcV�^��!�^GګM��e�`[676��Ƴ7<���]��c��N�D7��o�,U�h(2����������;��٥��K��f���	�d���:�h�)��VpQ������LܻG�
���H!��>fDp�("R�k����!e}n�f��!`sAM�?�C��h�b��<q*�;� 7%F��[���a,�rzD8��V�mI�?�z��8'�l<����X��ࢸ	�G ��OZ&ٕ$�s.=��R~��B,~8`"�,����UV��d��<�~Ƭ	�h�A�@ǨG
ϔ6��s�\�TA s"�~DyffЯ��4P�8Ѝ=�P�9�7�%ų5&�6�	�� ,"����
F�Ǫe��@��D�� � :��|�Ea��	lbQ��g�jۀ�{�w�� m�����sa}S֦9��Fc�v<��ӠK�^<GI���2��/��$�A�����$��+H
�}���v�5Kk������^����7W�52��GD���j��KP/��6����ܹ�-ۇǤ2 J���C43�H�h-�����O��88�aπι$1���Ȑ!
Qq���I�!#��l��f6���s�Ka����c��v�|�x�(��\����ـ+ݜ��gh���]yvkU~���3i!��J�yA��C�t(+���B��n�r�,X�_tDn|�0����:�9��:o:��BYҹ�h�X�t��'L��xhr��o}|�Q���_QN{]�p� �˿{��6�)����hz��n�B�Q0e���U��ދw�@!��H\(���Mm�Y$�|�^9(�?ޓ2���O&C�v�H>��M��߉��ěI����3��	I]S�Vr�C�|Lrp@^��r�[��D��vt����'���N0�jQ~緾!W�nJ_':Q�ЈQI�<����m�����,&[���r"�JU��"��&G�iHv$�4�H�BD�S̙RG�K�bN�-������חWI�G�	�m�ޣ=�}�m�;8���{j\�2T� m%$�H�ґ�H	 ��4�xFF�[����R�(}N�v����� dN�H2�L�����ԉ�D*��Kg�KFc29%|
X�U����Y1Al6�t�B_���{H=Á��x�h�QF�U`iX�>AO��E'*�L����Q.�K�����X�rs�s��l�pV��@7��:N��(2
d�r� �cu$���U�����W/���F۰�n��Oش�+K��/�^�v��x�6*�]�e8����ի
6��v{��e�ՐUl�*�I��Ό�ɋdI�U@�Ӊ�ߙn`C��㡬�.�q�� ��6�#�U��΂��ˍ�z��\�o4�n!r�Wr���})�ݱ���&�Ho'dl�!��*�^�@�+W�͢��˵�@ի뛛r�R$v	��)�&%�1���>�b�
� ���g6\ϩ�_��[$��FV\z
8�;�\Cq�0�k̖�yɁ�=]e����n�Kj���p�u���=�4��cו����WrIv���-���l$+1�8۠R���-�6�똌�� �$�'��G}M %tI���,��1.�N,g:����Q<|I�i���饗�!�ɹ~e�EM�>�RT�-d;[W��n��E ̢��)�`�u�Ч��.4x�9�s�7L�D��d���#x:��t��'ܣ��v��t�t�>`���߹}_Nz��Ψ� �P���˼��9nV-�Y�����=�hP���$:'I��EI���=_�֌!�yj�]��I,�٣ǎ8a4ۊ�G�7������x_�]�p�
U�$ēOLAp��}V_p�{�5}f���y�º����jso���=9<�(��''��^�Y���ܹ7�k�E��=F�&Gg�7t�+P�1c��j�$>�����i_���fIa|ki��o��'�j���b_��ܴԆ����lb��|/���[�Kmx�00!����2M"r]'�q�H:w�<� ��B���u�T'v�6�������WK��=��l�p�ar�^�F��@e�#�ʴr�x�8��3!�FE@��(�)�M~���c���j9F�(�i�,��&�{RB�(*JW�X�p4�K�ė{��F��takK�.n*��P�c�^�pԑ��9Vﭤ��jk�@MثH7B'�/x��d�QIx�8j
����vn�~�d*��`\*Bp^h��H�@��i��s֕��C�����z��u�cݴ?Q�xW��kA���YK"�J�E��G��`�M2��~m�<�[�J�	��b'�n��}X3�?�L��yE�Gqo��W'��4�E]�pQ��T��5���v,f���kL�����S�	�$Fl��� )2H#��yѬ�1=57 fEP:tC1
�W��'�󌷈�9�t��}t`
��CM�4��kӰ7aʪ<���ѡ|��w�"��ZA�u#x:�쓟 =���=
F�2SJp�mFD��MqѴKP��9{����r���<��K:���E����f(�rˁ֢,�^��Ww|(._$w�7��	[	�RU���fC��'
�栱2t& x#�
�d\�vhN�h����ZU׀z���2�@��	p���m
�s��� ��DvL ��R��+� ��=��`��Dv�>���~����YB4�&��óSVz� ��RP|xx,>$uՈ�,)�j�[�m]�(G���{���Tǣޠ=���%��?��*�klI
�hp(Q0�b\0u��ُ��E��"Sp6|���a�X�j���Iƽ"j�H�Y�	�\���@��lk�U;?���ԣ�J�*���L�E��؁T�f��'�H�y����C� Q`���EG+8$\���б�64�C�@05�2S����[�OD�#FC"f�e6f��X�X�@i����$����ШK�feY����
+���Q�9G��9F������e}��	RC����&���ۗ�U��nHGA���)�͝����sA�J�����z;�;v����E�Ϋ���!u�G���|�Ih�M��}�m�1��a��.2��AI�%�(���N"�s��r͞z$:�	g_{�v�Ker�����=�d�bL!B�v�tBp:}�~iC>����ܗ��)�:����txBsYൕ����_�7^}Y�စ|���������o�)��՚>���I{9�{yQ��(�Zᩛ�O><_��Du�r��dUϻ��p�]CC�sػ!�� P��p�d&�/)�`�8+�&bz�5
m�r4[��k�ō�
�nQy�U�?�(�Q`��_�.�>,��v��X����}N�z�#�k�.��J8�jw��� �|��tN�r��~�(n���K^K�v����F���F�\c5��';ޕӟ�͍csk����~G�CS>�������RC��h���+-�N���],뒯�$׌}�&^YC_ǆG�5�!�*�	�h�~��UF&w����ES����-y��w�}���(��)΁c�d�n�^�,As����(��>���s琖�qE�'��cCxN�Ǳd@�Ռ%�1�2�̣�8Ȝ�F�O`�%-���YW�^��ɱm�+�yRy��A��~��$��3�q�8�O� �(�:ss	�1ċc
�� {E����\���٣�� ��щL�рW���wz�yM�B>�2�u5�#���Z�n i��e����\�uw�o�\��S�$<�53���`c�
4��4l�p�Nu�!�0�܄<��������\Ǘ/]'㽠��x"+�:��{
�67/s�=>:"7QDO�z�c�|�=r�r9>���b�1�ז��6�qxx$�Q���j@Ϊ@�"����xB���֪ܹ�	��e]'����:99&=�^�s\A������=9<8�`霤�(�]YemЦ@�`������p�F����eV6C����X�jOO�R�:��g�������* ���loo+X�������C�����hg�đc��������ڮ�-�d[d�����7Ы�4}�v�y�����UJ��b��EA�/m���{����:{��qa|�R��l�YJ�$k:�7�y�r�	�K�<��dT�&��\��5�]*���g�Q&�sX7�αx���� n���[�Hp���
N��e���D��w8�Q��t�B/�7n�|ޗ��yc~�VVu>O4@#�!��y\ ��������L)��g��v<���t�yN�b��Gh]��eeB����e�	��!���ټ������@%��´	���.&ph����^hB���K�@�����R�:O��={�
��AM�u)ך���n�^K���^�ӳ3�lD�� �~ѝ��F�g�����dV�$���	#�
A4�������u��' �3@1{�Zvl�GD�G�T�ㅇ����r]5No�
H���V��f��)	��&�e�MEĨ��B|�hW�tÎk+N�ӯ.*�s�!�Cʯ���@�	�:O��KA��9������$����ff02�ѱEL�>�j�,�.HU�6T������l����,J4��J�rU��IJ ��%6TTl"y�L����k,l���0 G��"BB�����P�z.��A��b�� {�20����X�-qcG'�Ճ<��M`Bt�NJ9k3E���9���2��7����L���fY4�}.��{����A'">O�[��)�1Z�*{��0�S
+�Ӑ Ƨ�"�'̥'D����sz\��UQ������: �b� �8#D�&5�@Ã�{m�#��v���� Y������T4�����@���p�]�QSS�
�\�F��"�i{���1ˌ�P�7rԂ���ɂ��~ؗ��)�� >��a.�h|��Y��*��#�1 g��$��-@](��n
x֘�(��^i�%֍��87"�,(Q���Zt�q��NMH��½����iL����/U��!���9i�������]�*ب'��@�O��=Fz�Q_���9W�����[V������r��P���U\UЏ,EI�@�Y�4��:ev�$)�z��"L�(�����{��urMV��z�gh9��c����<�j�U�2\��iK�{�w�C�� `*&#�#�jb�����p�WeV)�S��踺��'k��E���էe���M��.S���Ӟ\����K*g�?�&Q��ٚD��q�NXDYj�X�$����}�wus��Gw<c��D�JO'�:Qpnȣֱ�x���3T��r|�Hj��`�&�3f	���C�m�t�!��"d/%�H��@QEg�UiYq�r&">sm}Q�m1�=�<��
Q2�&�F [<�`�9�5j�0�T�s��[�~��<�8�'l�E���_��9�pt]�(���8����l��ϲ�~��m������xKK
c�Tۊ�~ʌf�m�|_2L�����G��GEׁ'&��u�����E����6e�Tp[\-6E*��3F���E�d��g:��w�&<2J0i���S�Ě�[���k��s���E�jl���ECJcſv�s����AY �qt+z3;� ��oϛ����yR�]Jt�0��D�}�H���5�$t�E�H�F�%)���"Y��[
�h:8Oo*�t@�I�a5�#�ݑ���4�&�<���vYy�h �ʁ~_'q�ޒݨ�ɀ�١�H���UFĐ$�Ȣ�(.*�xo��a�!�б���8 C��r�BC3 _&`d ^���NC>���L`����Ǚh&&QHz�.��%Z�~Zm컞��;���|J4������y�*�ܿ�Fb���>+G1L�XE#@8��f!%	�k_�����XHD����'� �ƤR���l ���y�,�����t �v�r+��%b4!��7B!^� "x� pC���R#��"�a�[�,���bD��_�����9�H��~cuC�p���"���u ?�R�I^A���0F*g�!� �c�hB���~v� �Lǥ���r��Xp	�dA����.l]b���je�<3��p�ڭ��7�x��������q����B��N�~�X��t̱-����-����x�
)Q7��;�����ёUء���s��e9ұO��&�� �Dd��'���BΓ�_��GVK�.���8�<�,n+�)>��|!�s�c��AMǮ����'<���O����H j+(�� Ot�P5�������W9��&��٧�,��/0���x¦w��53x���"�ah=�uM�������8Wos!o�hŝ����-�E�Ȃ~��/�@ϗ�Zٸt:G����}mI��0(�ƃ�af�c+p�!��&���V,j
��yH8�qz��i$0:�i;�R����F�E�!�ݨ?�|NEm��:&��B��8b�����I�qC�����?����O���l��2�w,�|��aR�d�$:K����fv��
��&�T߂lTj�I�B+ؗ�S?�s'&PDz����R�!��L����i��T*��h�d�R���x��.�_��d��\��O���e�K�:6��H%�Kd\��v��*-���K��)�8p����%-@ዙkN.7����#Oo�v�I��}[x%�.���p{�;����5|�Ipt�7h}�i\L�w2��G'���sC[.��4�<+�Ž?B�?�t�v ��
B���ZQ���d�R� ����H��nJn	��L?�旎��{O�������
e�{��X��8Z�M]����R6��������p�3���$X�|]������{��������prV�0y���و��i�����kt�3 �I��++��G2:~�t4���F�ª��~��[r�٫�_��,/�Y��A�7����� ��J/�`�.��O�n��|��4 K	b�\[YjH�zUǵ7э>&������L�5v��t{�R���kWm������Wi�6�:1a��7��4�D����k�+�� 5�==a����a������F�wm:z� ��qHa��`(�J��g���T���ƚ�:7p�Pg9Yj.Yg�+��G�ܼ��%R�����H�WK�(@W�4
��;���o�p�q���l�}%uF�	I���D�i�ў�?h��J[�z? �h#MY8������!�D�f���*�8(uR�q#BkE�]+�)b�1���yp�YD��I��s�f�6�MX�r�w�d����uXc�v��#dV+���
dN��]���"'hPN�=�3
v�#}U�]� S����HΉk�IV�Eo .?/I'�\nέO��=Y���~9`�l��.��x& ��w�z����ȅ�"����`?����J`�s��xH��O�L7�<�+��\��e� a�3����&T���O-��E�sEvN�Q�x�X����T��g���3�gJ�9g�ҽ!�ş��Iߟ�>�J��I4�����:��O0I��d�A����B����K�st����Zf��t.W��(�~�o�';�Pڗ.˃Î�U螮ɬ,�N���}Y���V��Ws�Pc��T�s5�S6�y�(���p�o��77eo�-��S�u
j�����f���M�\��aE�C`��'���_�j3{����;����r|r�J�%UЏ6�'�ac�z��lnmJE�%6�3��s��qdA$�KBGqt�:kO��YYD�la�kA�.2H��)�6����hR�4K��T�!�p#�8��2ʓKYo䑫 �R^�$����g"R�i�*,���D邌3�]M��EZ�����x��f��S��f-�h��ؘH��Y0V��y{��wh�����Y�ۂ�&���w�s�8����Ӽl�DH���-�����a�H&�A�]./���u��g�]��|���\�&�v�:�PU�jRő�ņ��v�b�<���Г��Tn߽k��Q5zǇ�����I�U�"��}�u��
Q%F����j�`��H���,*�A$Q=�j�N�R4qZx<eD?�&ttx��~7՝�G�Ȁy@����}*Bׇ �˄�Z��p�x���c�%^��&8t��|�1%nPR�������LQ5���T�x:������4��M{c�^���1�8#ϩU+K������ˁt�AD~��Ra�4봻�h��Jx�&Ќ�z/# n���p�9Q�*Cu�OO�zs��3�d{ b�*��'.؍E���E�*�y�(<{Pa��_(���J
�!}��&�5��dx2�
�B�����7;����EG�
n$g�g�"Y�����d�S�l����s?q����g��3c����FR��%5�=O���\rm�;nx�wͿ/�3��e!|�X�����ZvH���Φ�����������. >g�]d����3���,ʣ:���/|�\��.M]?%�g�Fh�Ȋ�^���r��K\n�s���
�ȕ�%9��w>��] 8�_Ԩ�a(&�7��aM��W|��ɱ^���?9���Ӟ����yB5�P$h���킻�V5H5�v:�ܯ矁1�X�����X\��ڦt����(T�F�,uk@�l�@����
��ׇ��u%��'��M#��ɴ�KT#Ͻ�@��s~Ez��ǒ��2�[PL�����_��<πr�^��I�02C�Ͻ�	�7V���~��gl!6�'6����5 ��t(#5�EAX�^�"�`�{�#(I����3aL<G�>�TJ�@���F���5�$���s�,�̑pI)�8']S���~�ُ���=�ѧ�t�Ep,r�?�n��{�G��E������1Z0M�cDv�@D�ع' o�-/��y�v��鏎�R2]��n�~PR�0����N���K��-�H0�+e��e����s��X8'袠;}	��f�a+j�6�

�H�)`e��k��d�Г��"�/ =��K���X`wD�\'���T��,�u �A<�#R2�$���3��*l�~Y=]-@��
7�c�7)+�ȱ��1��)�QTD�Pā(-"o�h�d�}n0x~=D��N���;��"U@7�Ih�s:<c4���������V�t��ء��s 
-�/�����o��h�M"�s��XG�,��x��ͪ'��Ӛ�Ι�*m	I��q��a&��OY!�S~�r��$i�1d��������G���b8t�PCP��N��5�r��y��2,SV[��ǁ*j��Sk �[m��m|�q�A�yP�ڻ�84�,t-�|�v�3p杳�ɷf�Ҿ�^��.����g3'�"���a�4����ϥ?g���	lDn��ߎ�����DB)�:��y��KYe�O9�1��y��1��>���^z���m��[��v��m
>�&޺-�Oo��DmP}�����[���Y��^}Y~�7^��+����Zo�z��y��r�`��\�>|ۑQ@K��Fѭ;we�|��������J�s2��	��������~���3u w�}��m"$y
���/^��,��`�X���~r6`�-�/�\;���/�V��LSq�d���a��C��[;���sp ������>A�-�b�^���t�0��? H ����nI��G7e*3��D<v�EJY��@�{�_�&X�q��	�=�U���E�4?���L�4�.\u�c�0B��110Gq`�:@�%I�Y N=�f;� 	(��$�D��I
��B��I/-��p�����\�$����=$����������,8\�l��3��|Wr����t�	Ö]S�gX^�������x�Q�Y�)GD���P��>A��^z�9Yi7�"A�3@��cF~�$�>v��EB ����
gu$��9y�㛔� ���
l���9R �/#�居��)��Sp�T�HI"�x&�A(�Bz���je
Ut|��<�i<1��s|�Y���8��F�����@F������K�� α�j�DF��)g�9�<z����:' �Y���1��(m�.p�P�V�ɬ�`�4O��9Zjac-����'ԋVP,Wٮ�C�L�O�i]�[C���R<�;�2 
R�E�:(�
AP� &Rfh�GTh�����U�Y��qø�_��?��� =F(��!K� � }���l��j��.�)
y�� ���kĎM=o���-["�"��9'r�I�
�.�nk�QD@3d� ����UBW��,�qީ�w��A�'��=<e&�z�79��ı���g���̗dp�)�D�]���s�x>��p��ٴ4Ɨ�c/��7-�10�
v?Q!�=>^0��w1j��ݷ7����Al�]<��?����.  O��g9�L���QD���_$}��k`��Z\��.�8ҵ\��ڴ��9����ɿ��7HoF�'r������e�~,�';Rl.[q\XT;���*`��;�ʋ�]�ۏ��-b�B�ʞx${�ڐۊ�u-NN���h�����{����N8ed�{"�gj�Y�K�R�^�N���ǲ�0vd��Η�:��J)s�q��q�4��u��.ڋ��Wt�'#}������%}5|�#5�STB"�)z̦NS��n֒PQ��Ve�{Kr�y�9:ϩL�,�et��;��c�O?67��~����&�&.J��4f�1N욱�s��3#�Fbil�C�����N� ���2O$(P^��T���E��~{è��$�y������)���d)O,r�J��wƎ`x��$�Nx�`/E�/�8�	�'��Q�4u!��.���jz���Q���]8�&"��癴s�Q�4L�O��X�+�q�H6��r;�{/Rw�%�2rJ����q佸��&��f:_20s
��_�0R��M��@et2���}Y]���zKڵ�4)���:�zCJ�79�b��;�ģ.!6�4uG���!T�\�z����0�I�Oz:$&�C��X=�B���SϚ�����{���u�j�h���0@<�?�"xE ��+z��fyn�}W��D�h�8�P�Ѩ�9�M(�#��p1_z�{�9R�rE�?�_���ښۚu�P�RN9�$Ya���Q��Z}V"�PR ������D}r�Zm8�#P�'���:�39Ӎf��➜I���knNg:oWx/�,�ɫ}B�^�����#>�������h��0�bv`�< lc�X5~��]9�?`��gÉ+�/�Pj�e2B�#l��^z\q���b�R�����cv�E��y}���ȁt�h�Z��k��/.p^�3�hj+ �| `�z�^�"i�[A���=��.b����s��Ĥ���@l��%��_ñ���3-�.�6�%��[��x���lp��q�OGM�d���+�R_�����_J�J_O��F,�����Ld�e~7?���f�ef"��=
T����:��:��s $�3cwS��c��w4��>̈dl��DV4ED�����V�7Ek�rAN������@�XqeK����ୟQ����sR�V ������E9��~�cv�J-�U��+�D�c5�����W^�k�ś�6]��9�u����L�9R�7B�Q���8��JN�Eg0��;����ے[�(Ӂ�5}���Ү3�`䊙s��M�5W�q3@_߱.�{�
�w�BS�� �\ߪ7�ǆ�%)@������V7&�������s������e�F����b� �z���Z��(�R��^��ZΑ+�ga�'�R�+EJ��^���5ˢ��.�������ic�v���9g���������A���H��4�E��Co���.�����JW?�`�k�zv��2T\g?�(P�t��왨jf����&�� dh~������ ��&o�v}6^�s�ͣ5C�sn�֮1>�a"���Z�C��x^�S;ђ{�i���}Y�d�u�>C�w�;4�#�&e�4#˖;�# 
�A	�AB yȃ����`y	�<H~1�MY�<J%��lv��y�CUݚ�L�k��;u�ؤ<<�%E4�T�9߰���^{�0�������}OY��{� ��A�ck�������X�]-Tò7vh�.��0"ψ2��Y�H�Y'�:��Yc�\���I���{sȡР�F�
���D�g#>
l���D�����W/��v]�&�/��ݕ�`��q.���n�6\��!SO��w�}���^(���pأ*7�S�ܸ�f`�kv�{����Ci�]E!:-���<�Mv�@�cܶn.�I"�k�'��<�I��ԃg�χB��a�����g ��T45u��ZԹ$��g���C���z�ܽ�Pz
���z����'ù�]�:�YYD5��0�v�K)28��j���wl�r�|��5'�8<�-IBs�9��[oTd�B�
%�j�:&�/y��ϋ��ׅs,+�M�TY��)uqp��5j�:����J�
9���*C\�}%�������϶�s6��VU^,���=�+�5���ݧ�ϲ�t=tWX��l�:�����]z\�ib�S!]b���c@�Y'��e��#U鵬2���d���s�sS��L��6*k*2���[ks����=��s���	:�B��P����,G'�֓#��������?�٬�H�߇��$~�����]J���K�d��!�c�}&�(��(f�� w�]=>@o�L޿s_~p뾄�ɛ�P����6)4`�Y������Vm���f�a����i47���_�tɝ��_h�~���Y�)�]t�|�	��d��փ��ѭ��hcy��5n`�����;�ve��YC��$d�q����V-�W�K���-���2<`��OJY�0�T�.rr���*��V�q�㰞����o�>-��:n�a��!-��޾��Sl�q�|�XT ]��ʽAt���Ix�%�k��_ʨ��@=�Ha#��m��Vn|%n߳jj�ڇ���Fk;�Q#��������*�ܸ���P��+��׻:.�4��t �^��9#<���(kT����eb5��1�����ky,۝9@G�މ�@FC�������9�z����Oֳ�����Y��<2v�@��E+��7�Ñܹ����f!�dF�qH�#KѦE��ڎts�BO�n}��4�T/�-��l`�&Їc`V�<�|��0p�z���L�����rv��6�a��<�����H���1�j+Xj�o��M�Қ�� u�����O�#�[�(usi�A��Q���
B�ЧBɱS����<>�˵�&�����!S#�{,*��t6�^4��N]�:-O�j�w�I25�Q��(n���v���O=Nc�X��P`
�ӓ��L����d<��iʔ���,r��s+�Fx����
��RD���o��(�5.1ά��3g�?ŭg=�ƣ���+pc�/׮kձ3���g`kgɓ�s����9�H񜟫`��w�Ѐ��EhAA�b�?M1�zr,�A��� A�5�y��I��dς�XVKW/���4w!w��>4~F2w���2�XU!A�\�8�����+?��V�->��|��>�VT��"+Ar=�&��g�J�$�T�8�`R�j;9Z��*��=r��Ic�<�3}��Աޗ�_���,�Zn������?��?�!����U�^P��>@�\?��=b�7^��ŗ������`��6E�PQv++\�2����wg��a�|e0��J�N�}�L~r��\�T�jk�r��% c��y.�]��L��Oc�r6�f��m6�A�����9S�����m�y�B ��C��s�� H�s�0U�ώ&�l���z�����S'C�u1�kl��D���c�y��w/�b�yQzG��XT����,�]�އ��ʂ/��I����o��X�jW�ԧωIä�r�ڊ׿, �F-�(�y"��z=oh�Q�?��ɔo�c�@O� ����5+Հ��G��)�BJ�3�����uWCO4�a��Ov��{��E����5%`|�5_r��h��%<a�N�o��P�2�Bc���c$�ߗB��Ґ�nl���r���*�)��k�� �+��������])f}�y�\���� �u�3V]=Q����5�}��G�SP�$ݽ���M鏦�l��l)�62��ڗ���s���� ��p4t-��=Ir�iO��'�K�_����&�=<P����5)�R}�ƭx�pc���D��:�O�S��Q���t>)���Ð��ר��(+�kV�;Aם����G�!ӯ���j��!WFoV�"�3���QDP{@��y����<���78*��lS���7<f���NJ�w�5^�����Lfg:&�MLF���1ۧ�&3�����=}c^��F�}�)����h �T��V�ړ8�!�$ykKf�0�Yxa�O&��P�b͆����k����˵K,�`s%��Q)��
����m�򹱣���G,����w�Z�=ζ`��<}���\�v��`3�4�{.�(��(�3X>��2���/_�ו��>H9Z�J}�s�TA��՝^8�y�&��Jֻ�U�c��@T��A�����O�|^<�hc�.��U����aA�����a���ʫ�xhPG7&D�s��l�hh���zAN���o���7>�֓���ޖ/�|]~t�P>zz"�ֶ$���<��w��:n��2����ey��-BM�������4oEa��t�!;=~Zōft��,�;�P��g'�Ӆn������1Ԭ{N�@��ڈ4����RυmB ���&������^���ơ�
Ɍ�Hf�ޗѬ_\�|����o`�#�Q��*e�,�L2_�ɉ���;�����GksS�<��{7�AjH��O.Z;�,�dR-ޣD�3��C�n�o(ؘ��9	��y)�Į�@���k�j)J�2��Zn��ǳ�B��{���ٜO��(ц��!�>"���50��>d�*2n��S�L�f�lBk��2F^�-�4�Rs�[o��b2�C ����*E�)iqPн�ۀ��|�?!��]�������ZliV���U8boa�OFVl��n���%M�ןWf,�TbH���8 �{�)Ճ��~p�g�5�ڪ�ce�k���2"_����X�|Q:�$�k�h�[���-<5F  Gg}�!�T�����O��|�m��?���?�F�KIT౅f-6?��#J����v1)��	���p,�ߺ���.�Å��R�~]i6�A71�
b�2f�!����O qu�=��oM��������v�&g�#Q�I�7.چ�5laa_FUu�ġg�P�@m��"�߸/������y�T*��X+){��QjJ�(8mv�.zh͆r|6���L6�ޢ�}��y��1-H�4��E���D� 7�
�j��ا�L~��u9TP���,��`^ �I���е��~DAaԥ��i"7�Jp�`!W.�SRg8RԷ�N����'�n�u웱�����޵r�ɑd��p�hƐ�A+��=^s:�3�@��V�F�/9z���,b1ZT*[K�hښޝ�9�����b�<��J�^���uA&���e/����ZD����,�H���V�ԗ����5��`>�x����}կ������,���{���"�98��e�l��y�W�TJ���Y�
;W3 �{��m�#MǽO��Rq���Eǔ'��Y
�jI��؃J��]_���^W�~�C�k�jظ��O:���V	�S�c�/PI�v$�b�e�j��5]p�*!�=��|��@B� _z���`�@���XsJ���-
*g��?���ƽ�����_����	x�`_��Ͻ*�%�8��<H�&�_Y�3�����IOn�ۓ�Mi�Xmv���ا��A	8�6���:��=�ɓ�3�)d��9a-��[�AZ��V7�9m�Nu\v�3�>��Y���q�PVA��H�Ur�I�O��3}iO�Ӟ��_�p.z�Y�������^���l��xttT<{�T�ޑږ^���7ȍg��u�q0�Ff�\41/L��c�欹���� �9`����]��D^�]��M�06�zK�!�L�E���%&}�U�"މ[����-��m�O{����g>X��]�F&v'�3�ֻ��uw ���v���X�7ZrK|��G׊ǈ�Z��.1jXz�|N�Y�4Zme�2�[�@z�r��60�Ԁ�5v���?��r�GX^KXT�u%
R�C�2��٘�q�V��Ո'"���8ξ�e'�.�1E+2|�H0��9������z���1�|*��^-V�'�]p&��G��u�[K8��u 2�'��ԭ�'��7	�67������0A7 �{��ԭ-V��:f��Sq��cy�Jo�* ��t7u&�4`ڐKa#�7�����<�#�����%��s�l~�����W���Wep�Xv:��3hp��E$퐣�cb��k�W;�ᝇ�o��QO�
S���{D�0,�9;P����&��7�y�#u2�_��ȉ�/����^��;��5Gհ�q����j�!��@i����;w���\��P3��x��V��y�,폌J�f��3���E�2��<<>��<{����-���>�������ِ�iP�l"����E�q���w&?y�����pЕ��7�_�[���nw�qz'v2��2K�<9ǆ)����w=���r���H,�����a-�
����biw�5`��Q���[0	�o)�8��K��y�ꁴ�M6~�Z�����ޱ�Cf9��|W3��+İ�'���"�M�24�5�j)����`%u��[Q��W2f��x�,Y1.v�\K)UC	�d��֊'Ж�i��W��������n~,��ר������rnXw��W��$P����9��R�+���X;;ڄ�Y���)�`�%����>�����ˆ:T��q�x	mA`s_��ێg9�tQ�ݿ'��艼��&��K_���Mu�����A�IU�Ic������Bp��L�:�J����gO��6r��ɐ���8��8n89�~j_=�VE��h����Z7�ٸն���7}�]Y�EY��VK���y!��g�t�H^;�+m�������t�{�H-�7tn�j$������:����{߼q�'r��E�OO��ȳI.�Ʀ�`��შ�a�p�yha�<t �X'`^联���To:j[@8k%�y�61	���{ah)V���(�����u<)D�����k����M�}Xv�)ϰ�1Ք�#{'�./�a��^�`��p��K^��ƍi]F#��׏6?6$�Y=��R�qeWA��o�0QY7��<���*�N��u��y�E�L�c�\�+��}�q��XX7<��U�d3��:�|P��]䫰-*����y`}�sE�L={�
FK��/�
$)�`�P5���`El��{u��3���\��|$���H_�H�s���lퟓ��L�	���2�s�'
�c�Y�sN�{����ܸ�D�(N����'���hK�<$�Y��8�ػ��ZF8���G��S��ׯȯ����ۗ��?@� v?(�v�>�
��Yz� �|��ʭ�}Y�6զ�|5�*��x�"j#�Á���t���g��1K�28z$޾-���/��W�����g��ϓ��) " hc�M�9��ۖ�Y"�ޓ���?��nܕY�����q��Ǧ1�?�*}���m�͒����v0h�����yGל#y��X���g��]��_���)��^�:�^ �(�O�rO���;��]=t��Aj_�B?ər�e� �"ۈ��vr������$yͳ���n=�t���2�z[ŜE�
�1b��mPJ~4�s@�
-r�nT."�N�Y�4��ϵ�.��BRIo♨F�N�D�n�!�V���^�V"�Y�
���� z����X{�j!E��T���� �;�����g��XT#���LKV��?u���W��ED�ъW�U9.{�dU>lM�����R-&�q�$�T����*Э�x�.�V#Yf�����G���zB%�t}:U����pE��s�xԗ���;���Kj7����uN9/)T:M�ɡF�#R�Y�r���DAډ�҉c������S���_}�2�$j���:Ef�2lid�[��4�����Xf��8���;��Уn�{{6�S�*P#�a��VӉ��'�6�NC�t8������M	Q4��!z������C�c�Oո���Da�"���C�L����r�M�ɳ�7[��77����Sv�E�?@䑓��H���vx(<>���=��\�xs���1�#�.ԳN��GX�@�CQ��T;�M��c<P/ HgP=�:���^�">iVFi������\K�=)3��:�u��T6���^�U������w�YV!�uD�شW��Ȍ��oy�Z�[�WS�>�U,�Z �Z�^��m�t�:��X��HC�Ѹ��_~n��%����0� �x��<e�{��	�j�ܳ/��Q��z��Y��j�l���s�z�?bF���n(�p�Z8R!�n�d�N��s֝�&
���|�e*��a0�8 R_�+pY]_K�&g���4\��E�F���ԥ�Y��|�!A��릂�'�˽�wt�~^���ϫ�ŔI��!S�ͺ����*�;|t(�'ߕ��ߔa��"Z@!-�s� z��zͲ,�f-y��ꂣ�'�S�� 7Q=g�;w?�~�T���o��ξ��vu�f�i`�S׊t8����?�]�%}=�76������m�ӁԊ��r�;9�?v�QFն��%���#�<�fz@\���yO���_����mH�U�����(�n�M;U{���cy���	2��Ϋ�փgC�A���E ���7�I���H?�o���_�\s�/�A&��p"���L�����Wes��۴�S}zj�����rSA����r<8��֮G3�'��m��e�0�u�t�FG��Xl5����&�3w�����#���n��ɂ���s��e�]δ6_X��P#�M�Zc.;%�&� 
�������!U}�YR:��6MF����m-t�U;s�eVq&WSզ��Fditq��\>D��ԣ\ڻ��\��r�zp����^s����FQj럣�9�-m�It��x�Z�X,D*!��L�+��ΉgV��|�Ov$�J�W��k��Fg� ��%���u�%Ɣ�����8h0���<?�V����&N-������M��������H���|�O��ժKg���v�V�� PP�L�y1K8����/5Ag�.�l���꼶$����ؑh2��k,��--���>�C�>}�X'�=��:��-,�Rvj� GZ$�,��Wm3l�uu89�H�h�ڔ�vG�z/Wv��7�]ks������=x���F��n;&��CD��&��U'�L�}y���.V.������1��S韞��*� ���/T�b�'gcy�����;�ʃqBBeC:St.���d��U;����H	�1D;H�A9��#���B��'R�lE��&�.��ϯ�WC�57J��e�=��છa���b��.���FG$F�c�[��Q�z�5Y�hhC���O+�7��a�C�* �����1O<XX��%g)В���t���:��[=�����v�z"e�kbo���q�,7~j�Em�9�@�=��s}��6W�:L)�n5e2�1�1�@�i�,���0�gQ�����x �X�x��?�O+lYu'��(����y$��+ �8d�dy��'b�_gs{oAd�Nw}P�'��]��	�#�������W2RѸ&��<�zq����U��S��sǅjP���kqm�:�Zj,#��
g�O�Yj��˒�gW�������tO�C)�9��SF��~����fy�`��|���W��%���5�r�h=��y����ɩ��Sy��G�ß�'Gh����u��.�yQ#�Մ�����^�ŠAc�1ս�*��p5�0H'vk�E �f,�ͦ�Ѧ����[ߑ��c��/���s2T�	{}@�u��Gt��m�~��~З<�H�C4����a��`�O?;7o]V0_Ef���%_8/j���[j�&2�H-�- ��T�?}$���������W���r����V�'e��t����_��ܺ��R;躂hnM�o�M� ���}�e����zXw45��6�_z��pLt��>�k�
J���T~���ҹ�|�+r��vei49>�I��k����#�D
�������C:����mh����v��p<fy�s��0a�m^�q
Cr��ef�Z�X�سh		0�5�9"/�����L�R��9k�Ҟ�?���+���yB+�8�@�c5��K[��\?Ou{�W6i �&69���:�A�r�2��m&��\�?��m8Q>��6�-h�Ϧ�
Z8�����hX(�&�����G<&?��m�@��5R��9��eީ)�Lu{��!D��0@۪���A�����l���;�R\[��>��G�7�W���� Ύ���<�$���1ƽ�9�=|%:�zث��{�M3f|��#p�[���G\k>����5���5A��%�z�[�-�'���?:�98q���90Q�Y��זZ���%�=�A���w�v��X���Ea\y�[f���!��-,5��7�l�.s��tu Q�K_O�������sKIÆ�]
o6�c߰nU��"���Y�����ml�2�F,�1Jxe2�5� h�Z:�����u4��y��һyW5�x"Nhf���AvFR6?��#y�ܾ�����9�t5�B����H_�oZ��FS�ud�W��z�ґF�K��rJ)o����l�F5��dz*�Ӊ���L����-�|*�^zQ>ҟ���O���i�l�[�H��TatC���Y�ϥ2�(��I+��2�ZJUǪ.=:< ��k(�p)0�P���A������Τ��4.q=��i��a�t#L>.� �u�Q)G؍f1#9#:V0�=t���t�(Y@�1�;q�X��@h<��
D\�$�p�{��붛�	���P�נ1lp�k���M-�ǅ]��"'�:���遣zQi2rF���b=�L��N�x� T?���zx:Q�]y�~�� ��~�d8'�@BJ��Y�,c?L�ip0cs�ۡ�@~G��`��F:ɥ/.:�׍�r�ၴӣ�$��{al<��'
|��nl?��[iy�f6���3wΝc�p0H8�0��+�衅��l*Eo&�:xMf5�H�g�x��Јзu����l`��܎}�(�����{�P��-]�-�����!��5_� /\�PǗ�Nᳶ��*��%	�ߣqD�B��F����6v�d�^鬫s(��V/���r��M���pt�'�����^]���˫��o��h�P=�R�E��[ ��V��Z�c��/����u��;�x�x����Czh�UT`�v��1���?�%=5�I]_�[��c�z��t�*y�H1�q��L�9E��*���[�Q�����CWF�1g�f�9�����0R�P��*y6ԵP��g��|�K;��_�-
�w��L �3<�J� �z�.Sz��IX,�7v�A���Py���`Ȯ.���AS���m!�$��,0Ž&w����)v���� ��k>rR��й�c
�n?�΀(�xyF4H�������CAzO硤���p�E'9�������;��*��B� X��D�샱)8��P������Ҏ`C`[0�c�:�!B;�`���������=�{�S��C�	��l��	�2w�d6��2j 2# >q=�q���i��=��i�>��R�=���!o4.��I��,�TJ3�4-�4~mz�4�e�̃v�-�+�:�O����2*d�Ig�N?Q�Yf��p$(�9!a�`}������dϹ�����Ԯ:�UF�������ї�
�ª�|&F�� �h�	�H��8���²��l"Mұ��m���D��F�Q���om(�à��|��^U}&'��/���H�E
`��+L뫘�$��T�t��������vu��{�a�u��=x"C5��vG^��luw�`Ej8��'��Zp$A������̭Tۧj$m����������������_�-�@݃�A�z*�`���E��i����`	Ȗ:XV]�4^�z�g���Ū �3�|�`�a.^�H����#�0�'���&�Q��<�����r#��q`$
b�q�c���Pk9o��Ltk����q�K��j�t{��S=p���2����nX����7#Neś�d ����6�!�7媭�d٫��j�bs?bڸ�1G��E��hn�6�����n�qZ�q��f�A���c77�ȖrN��ވ���U�Ӡ"���8E�8G>�:��׉7*����1v�k4qXìf-�0ݚ�
D"k�� f������N���Qp؂���l6a�6	,<h�-B��ޔK�.H#K���v6Y��EH� |�E��Ty�0�GL��6vc΢�I����8`�g8��#�M����|�6!Q�_g���W�\��s�lX�9�߀��LR�H ��[��^�}�&�vF�a�@*ĨQ�ù�{�ŝ��:��e��<�\�P��%���<�cA?�����}�.�c'y��j��w6(#l���F��ў�&4u�Cg*n2@k^��ohgJ� �#��
�B�,�Pi�(l���T����k��OF]s����"E��:�"/mg�I��aM#�9C�^�bH-d/���ӇYiZK���'�f��)�|��(�k�D��I)��^7��p#��a{�Rx{�5�նFH1�F�"9��O�Bp�ӳ![�M����,�5A� �o��W�d2��@U-#�>���C'Z>Ň֥�� at����=A� H�{�l�c�fu���������tA��i���P��ok]�X���մN��}�Ϧ��{��c;��#���ԝ7p��䴍��#��{�й�u2�6t��8Q��N����5(����/?�7Ÿ����f�ng��o��o��8+�Q.�:ᅞ����q�-��
�`[q���c@�"[�l��5�3�a��Á�����sc�s�Su���[�����/�L����, Ȯ$9G�ae�*��E��.NӍ]�Й��a��X��wD�����:Fu ��� /�Ƣ&;_<ưT~��Q�v��˭N����Ly��npړ��]�W_�0"�v}P�FziQ4xЦ�H�w6e�?�	�H$P5,��� �R��#2�^!�nw�X.�+x�1����"�'�Ѣ�S\�!��<Ԩ��t�INd<<#�2<9!q�`�-��k_3a������V��xTA��y��<�0}����.S��qf�V��'��"���E�t@�]��S�^���wʃ�i��)�c�f�s�aoow���:����E)������],k�o���f��t��>�`�t�>#�d>�� �㍤�;��~���n)#Ϫ�2�hԢW諕=H�-��_���>mQ�i�Z�A�øV?����6�Y�k����$u���=]FE���#{�'a[ZF1��gj��Ƙ�#��p�1|��N�%w����y��������,�FP�Ծ�r֊-6x�L7ez�:��6��	�w�jYV/(a�Ul2�-�VQ���l����~���޻-�{}���H]d��Ҝ?��M�.��xt"c;��Ģ�h4����-���#=,
�r��kn�bFz����JЌ�	����>�Ă�������/R·�v ��scyJ��@H]Ǳ�����	#j����������CA!2tʅ���u!%��n�0@D�YіL' v{��hc)H�&L�Z��j�;Z�^$�#FWY��4!�3�ã�}�*hW7L� �#���g����Z����$3��C<S ���:ʧ<���Ђ��9O(Ԏ�oNM�Ԭ��_��LI1b�*"E(�!�[s������AG ����:��schY"Z�m�)�:s�D��͵�F�����"�Q ��I�/�Y�������A
]�C���]�.mg�j�3g���yde���>e�on)w��]��l��`L�)�&��ܥ��i�S����|M8����L��=R����$�j}�X�3:����$N���,�J�5�Gx�fӭ���[�dQF/�(��iv4�F=v�HF8�sA���} aFʖ9�ܣc����0���͹ƀ0?��Z�yB[���&"[�y�s�mqOw�+�J�<�2�S�- ��%�nZ�����9'N$�P܇}��b�Ĵ�<ܞ*U-��Ӌ� ה:�=�d�*7��`��o���ś�+��MuEl.����lk�k�9G�U�+�L������7�����7(�5�����R��zm�̏G���i����<�:�����ٕ��h�;�� ��v[�a����w�0�ݬ��[I���ѕC�ռ8��:��׹hu/롓��!��Ln\9�����v�U ��y7�L�	r< ����PꨌF��m�m�<Sc�L?��S.��Y������� ��x^� ��&]}�	 �I���*E35��A�E�	�|-4�tQn�b��JdK��L���@���qR����h�s���H.R��3�����<a������:�9�L�����N���\�!|�x͊U"2�A��Y:���iqx�	�3�O�%x����D�~�Y�cS�,f�r�a��U9	݌�g�Qe�8�����!s^�(���UT�ǚ�c+����uDÜ��Kn$c��OqPl�ϟs6Pa��0�&gj��j=�΄��81$�G��.����d���A�4�(�@�F��ٺ.4�=�����%CuX��~{'O���a��GM��/kR�� >��ߕ�}#d�a��ꈫ�c��(R���@4 �`�F5�D���Mu2�����c�OW_��)L�h.�=��f[e�bfIsa���Z�)�)*@��(��k��zv�T|�׾���r�����5gr'�q�9�ذg1S��	���1Ra	�CR��3+6����R�
0��<%I��<��inX��&eb���Zق�#P��{s��8� ���ĤI�P)B�*�A��uFR}a҆���k�l�l�WGm��T��+��eу9s�§�A`�Q{;� �k�gyY�����+{N)����8�{���s�2CRݧ�{dnb��oo�|��;����ק����������m�|U�oxO��+����9\����g�՟զ��jk�`[dk����+����~_����U�����7�?z��՟�����������<<�]]�]g����������?�����O(��ُ��=���J��    IEND�B`�PK
     ąnY���T0  T0  /   images/5107842f-df24-4ed4-8dc8-476b8a0f3ddf.png�PNG

   IHDR   d   ,   ��U  iCCPICC Profile  x�c``\���[�$����WR����~���A���A��21���1 ��'�v�.��b p��'�@�\PTt�.��;�):
����!�;	V�d� ��H�$$6�.`M6J�DvHriQ�)ħO2'�N����&`/(m��Qs����$7���ط�U��gլ��_{��K���KR+J@���@a�6��E_�' Ēf20loe`���SY��������< ��Mۋ�l�   	pHYs     ��  .�IDATx�U{	�dguݩ�^�U]]��>�Ͼ/�w			B,��cp�6���I����8��� �"!FHHHI3�H��=K��V�^����J$�Q���������{��ﳞ}���_���4��,��9Ӭ���xh`-�_�ל�H0d6���X���7���f;0M؆�@(�/K�Z�)Wj��J�0�,��` ^.Vlx<N8��7�Cm�S�#������ 8�<�'�/��
ŕ�?�U�U�k�L�qo��R��oo����E_�X��C-^Ӳ~5�cqM6oǿp�msU���;ar)�;:�2lh�=f�\�ةl>��~�l
���T2�[0=\�iڦi�Pu�fY��[m����-��w<Fb9���ۭ��l�Vj˰`p&�0�����*��Ǩ�z4�k(WkX�
��L�D��]��Y���#oM/bWKCi�ɚ�Z+��1�
�j�S��(e`�#0|@���%���8t��Ш�2_3`�l~��i���{�
���gm]�!��s�ّ�����IT�$����������P�V7��|�
%�j*NM?����'Ǳapm�� L/ZH��x��\��,�Y��U�\W'?�	j4�_\�\X\�����7�j5���%���+SvC+�Wڎ�W�}&/W����J�A��ܱ���Z�W�[��.a8�J���}C�?��ڻ=���'O}�o^���[)3X(��f����M��J��-"񡧳b�F�,X��R���RyL��XɔP�t�S_�G6 ���:��V���-�!ackgX��Y���i�Z݉�XG���$t���w�O�nH�0b�� ��D�����^�)3hM�V�:P����?$��6�*�v�M���t6���!��G�4�=٢��\s�f5��	�엎a�ܠc�0��(�}�ή׾�?��s��7���������wl+��~��_��B⡯������rxf�Ƃ �����F�2�v	���}�&��8���8\|�ZvaC�U�H���t��+�I�qi��/b:[��(��'���5�j|��q��l�WQ̗�I&�n^�bE�4+]Wh\sm��&�*�ɺ�5T*y�r�wvc�Z/���P=�<���[�MV:�#N絜*�4�ޮ8n����8�c!�LC?.`n���Hs��9�Z����8����F�p����,��G_zmq�?��ަ�u]X�f*d�Z5�ҹ���W/��B�
畿|��j�5�8��g�A<t��=q||�0v�$��2�����6N|>K�R"l�V�^/�6��M��}�x���:5�٢�P�J���xO����r� �td�^4�2����D��u���<�}��v��Z|�N��A�67�����:�׸��H>�w���D�2J��\�S�åd�"��A��ŋ��Cx��0�\]�''���:�A�����+�����]���w�N~��7���1�ڪex|��T�����f���ᇿ�O���Xq|>n�B���C���kGp��Awɵu]L�Q-YQ*W��ʕ��}0F(Rg��s�P@�L#���[G��������#�Z�_˨��e^��\�:W,o�\'�Y�X^�=�֬s꾱���@�D<�&��\��S����T	 ��q]w>}�f�b V��lrͽ��[�Ӏ?@*��5�F� 	(�!��Kp��߄k:��ç�����,�[����s�{>������ye���9��f��L��6�Z�^�,~�o��+�z�Q�4�0me�״����څ��F��� _�C؃,�ʕ�8u�4��8���d�9���:b �����o������0��Gs$�/߽[���;o�!EH��+�P�Xc#��gPcD6�\"�E�ƿ�Sw��v-��/����P��g�����{l���#�U&�5��nf��s=5��S�~g��{��8N�9��)`�Ik-��hkk���ضu3�7�i�OgstVܰ�����_�ѣW�^hƙBm$�F
�-���+�[��D��g$WP�&*�(����0����5�K��B��KC.0�Ȣh�������+ �%.��d�(��)������yO���غ}��G�qt�������L�/�|+R8y��?�	54`mu�lkN0��{<.�UcJ-gT���$��RX�I��!M��e�2�,'�{J	���ܴ�a;���rBg����L�y�W��/~��c��2!��\�NPܬ��8/�ka˖-x�}��k��Y3���������[�M��/��j�@�h y�"�zK˓w{E����� ���'�����_�� �lˋ��
/���|�p��qMs��p$�R���q��h����|���S'�������ޏZjyq�l��fJ����Q*�����k%�7��D�Zj�����@7.�KE�H�*�Ѳ&3W���I{�>�u�6DY��nX���$�bK����w�m�hM���fu�~��s��GO�P���B"X���l�ZE��h�#�Ǒ��Ƶ������SDz%�xc�|�����޹�r$�Z�`���}�&A�F
����R��ᨉ/ݳ[�vyq�t�ı��os���Z�d�%fH�?��Y�&q`��.�҈�а����8q�$����Ձ��EܺcKkY<��q|b	�4�P~C]m$^�c��F��RMG���S���{�F��rG#�إ����_�b�l�ct���q��?�ɇp��a4�d�������_������Ng`j�I������2;��`S
A��T+�OK"�|���=_��#��[��J#o�g�>�e"ĉs@�%AC��g�U���k�dq$�Gy��a�1,�ϫ�;������~�� B���q����81^�Hĉ�%��P��)����Π��i41ڣ��"�_���N���|�Ɲ819�'����A�}v��5 ����|~xEP9$�7�1���su���)�|m)�`"U@���#t�w�w���c�F����(�#�?�?����!��b�HօX[[Z���iT���)�&��>�����]�^�v	(�����+r������It7%�G�o��vI��r�J�	Xd)�0j^K� ���-m�is�Y���.�13����h�"�Fkk�[[�c�HQ���q�=��&��*Dc��_��*ic�eQL���k��������I���v��o~�L�e:e�����EF����Z&,�ɭ�)\լ _˨*�U=w��)��H��$�}��I��r�����V֓E^r�,�T/��2~��c.q��m-h�7soa��ⷬ� �k���������,�V]�]g|^f������[4%q�5��Ja_o;��؎��"�ZYb�"��X
U"���]���͢�+(�~�?@����%Ft�����j\)|%jqJ>�����$K+W#��CݝhN4abz�LmUcHz�����4>���"KU?�׍{�?��aءj�]��p��]��t*Xd=�x�K��~f,Ӝ��+%]�j_��
$W,v�M�w�>���������\�|�%,��%�F����C!�L�-U݂n�>~�&6�
��![��������2VS�Z�jwC���@"֨h��q��.|(��X,l^�m��Y�ngf��İ���E�ٟ���%��[���N㒉J�1T!~?i�d!Eޛ�}�.�	Gx�֝M##�4��[u�����^�5��έ�)4s��=8x��qm$l���;q��4*����<a�N��I*�=�ꪽ��%a�z����Z�\]�{o�!:��7���E����X���2�v�܊�xXa8�˹"W���6	k�$Et�H8�UH$vmۂ˓Ә��su��К63=�'�x
���g��e��ܢ���d���[��?���]���f��_�Z)�#l�F܀k@�B���S4UX3�dZd22��E�����������W& ��Ã�t�SӺ���g~��;v��kK`��^L�7"�ZAaq��AD��p����b�^r��I����B���7VSy�|U-� �Ͳ�{{�c����ݭ4f��؉J���O_7Ed�ڣ��X�H9'�*1I47���(}�j68d�����!*��e�"B^a����W��λ�it�����w�g���[���M�Td�`y�R>+����"�P[il�8�3is�|��a��l&O�Sv�#�
ɼLe�ZD���kO��kkiV�*M�1a"SWi�>�e7m�Cշ�צ��F(��ny��a���ɟ>����4�#�[�gt��,a�/�W���	�x��8&ג����׎c߾Qf?� u��"5�֮<�z`S?FGu��<�BHhllVDu.lL��:� <C�E�ah �^��>��ǐe �B��~�տ|���#����(ll�# ��h��1��c���6r��&��#�l�QĘ������3
eU�C3E2!
+C��YO%5����%֞�����q1Rs��6ҹ��~�� ��}��	�n�����+A(t�$�6܍�����-xZ���u��He��>:+@��>}����0�����=�qni'�Ҹu�����:������ɚQES,�TYjK���8��0nmm�>�)��xpAlܼMY�:�D�z��k�.i���z(�K{j�U�9E�p8�F�P�b1�02A�cG��.������Ջ�ή0���MQ���7A��SKOI0rb����N�)��)������WY��FV^��d��E�iS��Z>�׌���I�M�U�ahx�d�<����k�Iހ�mDk��F���5��U�w~j[v������%\<w6�j��A,k�>�N��`�؝�W�;�6�M-��ٰ�-�f���xc���f�v��_���Yc3�S�V	�B�������QH��T-�GU���J%�Q1X����U�E)֓��zx+nO�Nm4�@�����t���dp��_�%�(�q#��2#����&Y�������T��$SRe�i�f\�r	��Oq���
�Z+đy:Q�M��&*���EeX����W�e��4k�(do�ꚴON;z�o�@�j���'��ן�^�X?.ↁt���)Ȓd�qy�a�`���e6���$^8sq~n���}J�U�K��
ٞ�!Y3�|�VH�$�����!��/0&53�Lj�ʲ�K�zI $[:���8/GyE��x�KK��fk����I�ٱ6����F�
�r�`��6�)�,-,�BKF�'��Ӿw��+3"Z�Z��L�$�tӖ�X[]���"�MMX[#�"t����iT	�hok�F)��i�䆃!��F�<i}ȵ%c�桃�Wg�U��)���͑dh�\�YX^#��;���J���7����
�=<�D�Xb0	�=�������-���٨������?"�,�R[���i��%�z����'h� �]2BOE��G�"t��d��
��A~	l�ѭP4!�Ժ6 �;#����h؎�K�� ��æ,Q����zJWa�Nh�I�(�u�RĤvod�ـ�o֞QS�S��3
�3��4#M�l�����FJ3NT?�-��HدuJ
�'#�Oz&Ej�뙬=>:@��BBa1��X�Y��zx��LRDhj����Mz_=��C#C5��Aq���$�r�
aɂB����Q�6_B"�Z^kbvww�a�{>"Y��8�PKW���mzr���*�MQ�)�%�K�%�G,)�ҟi`D+W�F��乍:~�L��.�'.�<>�����¤$�qF�21����9�H4ɻ�Y$۔$�	d��2鴖�0�.Q����k�t+²]mW3\Ma���v�i.���n�'�j$=I �R�'���q`�v�����@ؒPX�Qғ��yS;�������p	���5̀`��2��C�Jg��UJ'â�B�mY�V�s����;l+a��z����Ś��)-J���8����dXBT�>1��prI��k����&S�I4pW�%�yjj>O%E�BV�StbYuL@��`�ԭ�ϧ�Z����[2, n��j�������P�Zܩ�q��m��Q����+�D��T���Z�ʟO�ױ-���9�#��N���	�����ݧ��D�������(7��4����(|�� '��0�y��,�?ifh�\%z�CyF{H�8D�'��hlԾ��(��j�hg���"��JF�{�}�Q���07?��@��{D��b�0ʂ�
��f��������
S��bZ)�22�msǨ���+rl�-��H=��{�ɼ{\(�YBbs7��TXY�/	C�\�Y�)���~�ҝn'�㶕�\��}�^��_XRc�c�8���&�°L�H����Y�zs5�Eܮ�eƅ49�evX�{z�I�/�)b5S*X=�R�������
NJ1�p���a(�I`�J'���Co�N�͕��:�af�E����q��Jc���h������U��ڝ����k�x�K*b����]?%�x\��S'5�u�j��P+��;u�i ɑk����=�i�xC��0��a���'D� r�آ�֓hC��Y%aYƞ�������.����19��Ò-�k���U�{��f�׻�9|��d���=�ٵ,r�JV�¢�W���#G���%nk玝x��׈���t:#!n�.cia'�������]���_��099�r��k�u]�S�
��V7��J�Di��{��D��h+2D����k�np�O�a�q�*F�0{�wn�����0ꇴ�Ϣ%��K4��t�F��v�ٍ�gN�C�B��Y\�,XX����3#�	�"	�d�謴4��$�l�ԺP`���h�ŧ39BRQLJ�d���0Z�Z��6��
��/�m����E���:���d&6����;v�@߆wJ!h떍L�=��ΞF�Q$�PÌO�낤.�n�9�d:�h�a|�*���gҿb��O0*�j��vaY�L�X4V�:f��"�[�]�ZpU��;�bו�D�i0:�"��YN}T�m�bvy��.�X�j����4�Z����o~��}�,�b8i���/�w�P��v����Ne��"|�-ɐ��I��nq ӌ����D�:Pŝw�FX�n?I.���P��ʙ���ZI1���2#1�т�����?|�{ګ�����@��,L��+�~	C##ڪ7�M
{t�<#���.����߫�D���TN����DͿ���i��iNfU\ZJ+�:�Yw>��X��j�^|Q�&|��+u��!����ϥ�U5��W��Ǧ��!5���]��u�vf?��2!�*3����8s�v�܅A���ܼ���n975�0�p[*fH��k'm���#��R&��4���?�*�1�`}��eLe+����*�Z��+���0
��j����z+�:r'N� CZS6"J<��I$!�N��ZPVA�J��dX�%�8��tP^+2CD\�4Na�`v�}�ضm+[B�)����3����(n�i�+=���rd0��:��G���,�;nR(�7���xf���#B'�plv۩�T�C���◾��{��5�Lx�42�GxJ�����������B����Cf��R��.!Ϛ�.�2	�O��'�iZ��/���TB�4���'|=S���i�lC��ّh`���P��ɟ|�տ֨�:>�ѡAȂ�����3s�9�W��s:��������� Es�X95=OV�UZ�u�f|��j�Rw��Z�`���Ӱ�k�$Z��!�z��S��67m׍]�k;;[0�ڈC3XX/�U�S�6������}�F�� ]'��Mѐ�a���ԧ>��~�;���h�1�rY���5��=O�9�@3� JV��">!۔(��yeb�fY[LBHʵ"z��8���|8�/N^©�ܻ���3��d�AC���ؽM�D��#t�Y�?�������7������7�ʬRI��<)xҗ��9��)!g�Y�?q��T�i:eMO�D��AM��(M� ��z���?�2~u�"�I����ʸ�!G����fܼ���f<��4.�{蜞�Ae`0���",Z�,!\H�+z����3�utQ���2���־n4%"�A���1����O�����.�M�a���mP%/��ZW�D_h�1��25�iy5U��r�{�a>�"3K���<���+�\Zl�*���̥�x����&̑�m��pU-�[�n��|�ﾍ��Y'�jiiAgW�N	Ey.Zg����5���B��x��yvv�E۝8ܼy_�3Z���!l�a=/�'x�U�]���ۃn:� � F�l��u&�:��Ȯ�r.;_�C=;>��=x��p�x9���Ё�f9�����2�eIw{~��5Hz,^���y|ঽ�'��2 e����PI�te��%6k�f�]u�ܽ��((����ɺ�^�t�F���a��������f�Oωx��7q!EA��ZEX�'��f�f��3�Ǳc���3�)���u����ٴe�����G�?��_�El�k�Z��m���|��sa�.j��ɩ�O5RT�y�������k+[��E���WYh+==(�.�wC+#��gvL����ũED�M�����,���n;�x^�훘�UP�6±<�u6u5� S��KHͯj����yl�I��1�a��+�x��9ܵ�6'K���0�Lz�����/0 ۘ-mJ^�+�cіS� ����1EA K�gk�=�!
��<��n�MOW�|��?>4����0m��y?=W��R�T ��ED����q�����H���ޖ/Tc$�)���G>�[o�	_xgΞgz�(�]][�ƣp)��|V=/؃��I6I\t�L��1�K̴���㘳"\���ujf�v⭫�:M"��ֶ���aN�ߑc:�ޜI�I�!62���wp�a��B��������{�d
����C��ٻ��-֊�g��1�{73�k
_7\�(�}�Y��W/�8��Ҧ������ޖ[�����o3���݁�?p?ڈ$�� Ɂ�`[�߿y�pO���5�����Lm�^/I+��wtjO�~x���kho�3�Mm3T�׻w����>t���3a];��8@cC����6n"]ܩ�^�z�Y��aV��<�/���6��,�~ݰ�v56p3bd^d68��h��G/��H3k�<sa*�
��t�H[3���WF�h
����=�Ҙ��wj~??~]��dv�����D���=�mC���ڍ����'�z��}�m���k���U�*s/��Hk��^���ܽ]��¾��k����1,��ea��!�D����-����+Wc���w�sS?�'_8=���{�������#��C��/�-�N
���>H-��*�M��P;�J��(���%�<V��2�������)<��j���3�=VNʸ~�o]�E �����Ս�ނ>��i�;�,�.⎛���ϼ���wJ=B��7��Bf���I�"!:���K���Z�����`��4n۽	��-ʦ�\����y�my=Q��I��Y=��a��G��Td�e�~��8��Ӄ.)��v�>#�jE��&��7GHb�Sd��ѫ~O>�T����CJ['�WI�h�3[���]�(�1Du����B�"��BNeR^�#�X&/�LY��i.�}h���_;��NLj���G��!2.�ƒ�����fE�'��Z
W/��``I����|'^<�z����ڲ���D�t7'�����_�#�\9�$��X\��Efj_��������
�?z	��9l�o!B40���?�����R#�~��%�:��B��&�85��8��s�Mc�� ��H&��2��.�A�����5���|��_�b��c�=���4�i�j�\ST�Ѡ���4y�ծd�N���J���*5B�����,|;T�r�@��Cxeb�u�ہ���V�9>�r�H�u�������a fRQ���&$|���(��Xd����刕�G�=vy59�H.N(��3�/��Y?��?��[�Kr Ĥ(ze���<��c�iiBc��-`蹌�	Ȁ��s���+	�Oyj�b��C��3��ёsH��%�a����Opz�"MF�\s�opۆ&�6�qy��7�S���
S^qpfq	_��$��;�k��b���!����{���ج��T�2MOKU�v}�ϝo
�`[��ǟzo,�0Q1�|A��Q�C�cC&��5li�`y|ՙ5x����LL�z��06�t`ª"S�Q�.�Ǯ�z�N,�a��ё�C<c \�`���0½�EZ`�����x�)�k8Ya����kwc��At6�!
p�r4q��.�K��ˣ6�����O"��#ZG�y��xn/]���]�X�N��x�n[���,'K5��T&w���C�pߎ�o���k�O����x��m[G0΂>��SM~륓�u�4��3�ͽ�h��UQ�����M�z��F��$}�r�lP�0C~{�*^y��_ZD�Yb��ڛ�n-�9�<��Q��}�v��u�~yvq#�ݝQ�޼F{?sj:���;{[���Y֚��/`��2���{n��SW1�;G�C�-�*h��,�&�i��RIO?x{��4�[�z�{��$(�)�2P(��U}�4C����A�1���
am!Yě��8Bq�Tq�Pn����+8Ƣ���q��Nܳ��/�����������f��5�E}O>w��#�������B�w��g'	Io_��`,ic�&�_���so�9�(����N�r�:',�Hf��.>W�"]ɑ�p��|aaS�f����X�!o7��g}Ժ5�Y���W�����E���Q�Y���6P]M6��t�K�a}yf���� ����:xr�h��0:<��s�(��b�q���2��l����!ы �h5[�SG�p�P���[:�Гh@����y����&��u�����ӬyGZ��~��F��-��|s�z�Ώ��/_y��x��ٿ�����+Kư嗩�:��-����K_)|�����5(�#`Ƀ.F�����m`�ѷxi�]���܇F*ۀ4��>Ŕf�L�#rp��<�J�u ϱ��vc�}8�q�?#��������(q׃�;O�A<ю���&l�g��Fa&vS��Q4�w��|�/i��$Y����ݿoL�`R�K���J(
�&����+��Ayƃ�|��i홉#r���#�²h�
�#V>/
^���8R���F�����ӫ8���q.=���K/���'>�}��˭%�?Usj''�~ﾽ�Ol�j?�黯y�?��o��IZ�5.��d��$��ݘwμ(�X%�Y����g����?�� �.1����LO}6�>`g�.���`4İu�v2� �$)_3J���R;6w���\�E���<U� �j�,�ѥ,�|0��i�G���&N�c�P�MD��U[�����j�����^}�s��O�Sm� �qɊN�K�z�!)#������D���$��ǵ�߻���\ǟ?��gv��=����e:��2��V,⟛�f�N^�5������6Z2��{��c�P�1�.6�GJu��=��?� MA�>�/jSf��_ϗu��u��ܸ�	��D,չ���b��D/7���t���]ݍ��#|7�ca:Y����"1|�!ʢ>��A,����k�m��mb�2�_%�WP����7�G(�g�%��}��fן�5��
���1�&�Ҳ�6赚��Ū]����˖Κ
_��r�Y&����=��P�:�@@�_i���
�+l��Z#a�����J�m�]h����_�\I��
�%    IEND�B`�PK
     ąnYP��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     ąnY$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     ąnY��ƌ  �  /   images/04d2d11f-9dbd-4a2c-b6c9-835d97151b37.png�PNG

   IHDR  �   �   @w��   sRGB ���   gAMA  ���a  PLTE�˸=�O��i�`j�Vb�SX�Ov�\o�Y��e�ǩz4+}:��l5�@L�H@�C��i��o��``b���jjjosk���fffvxvzi�������ċ�d�����������������������➰�s�����Z�j~��f�t$7(%8)RRRIII(O0XaFFF�ӻ:ZA:::000)k5BBB*,->>>LMM***" '''%$$=H'I\%Ne$Th)Zs(b�)x��m�.r�,v�.~�1��3��4{�1}�1��3��3��2$?*233888444YYY����pܓ   	pHYs  �  ��o�d  IDATx^�{�8@��6g2mӄ�� �l���4���yn�$m��>���Xݫ+��w'V|�ׯѕ.�X�lH(����`X��q� ���qJ�L�`�Y
g�0���3�d�Q�8����)�i�4Ə�BŽ��� .QP��@8CA�Z�p"ۇx��ju�ժ�K��a�=a�@͞��Z���N� B7��Z�Af�B�.S@ُ��@��~�VG/X�Ux�Z����P�7-wҙ�lG@[0?]�%;��_Kv���Z2ek�2[K���L�Zr��d�J��m�YK����YK�/TK���%ˍ�,�Nä<�*	P�B[����_D/(ɿ.,<��$�?]X�5��<��J򯋘�$�?ف�����g2[I�l%9O�\4+���"T�!����d��$�?YX|J��z&�B($�Vⅳl��fe%y�$�!B��aBK�����$���¼���I2f/��d��$�l����da��d�~�%�e����bc
ɸ1�M�evIKVO����O{%�a��GZrx��`�i��'��O�d�ʅ%%���s--.j�Kؼ�$�1|�%ˍJ��&�*[I�َ���Ir���
��,��J��&�fv�̶�p,,˱,%ÙOL�˅�ʲ�3vSi{�%��ZU�W1\2%�C��G2�K�dqH$KV"�*;&��aT2�͘�*l�[
ɲ�ޑ�
�qm}}Mj�],%c���Z�,[	�wIK�wD�s2X]�d�M��D6I�٫Z��&�*[M�xĬj�x@�l1A�8��d�V�1[l�$c�@KVO��U�-K%�X�Pcs=� ���N[66��:��B[u��S�z����b������l&ɐ-�NK�l�!1[,&��ʖ�œP��٢�h�ؓ��iQ��xH�:[IVٖJƱZ ����r �d\u���f����*�w���V"O�r� 0���`�A�J�S�)�(5�a4;�D���F�<�¥&@x0#x E���C��ց��D�2�`%C�M4�P�:	m�Kh��tϣ�Гt�=�%̖�E{�Σ��S$[:=E��yh����*-j��<̖έ_���fb���2� �P��#<S�]��Ӵ��K�:ۡl%=���
�&��l��HMZ#��t)��l�QJ�ҕT%]�ց}!V�=��t����Vס���:���S�%��7Z���� ��lQ�S$f:ۿ<���=��G}W����xD�-u,%땕 fd�8���d�̍�Z��j��^�f�E�V�<*n��٢�����f��y�A����pq�l�tK�Kyσ�$Q�1�q(�y؊���{k�sQ�,���P�\��Et� ��^E�\)�=-r��[�L��e8:xu.t{�WΚ8��X�U)Y_�8�I_+1VA����nue)%�>�%�u%c�>��n\�d����J�2�A@-��d�L#<���"|}�6�aJ�Y�s��i{o0�W������XUMJf)���7�$�L�����-���m��kP��ܗ�B��O����,�\����κ��7V����o����+yI�I~^�?�[��+�]�r�~�����-jpݗ�U�&oq@r��;�H.6ժ��oC�&^�N�bȑ\��w��ɑ̎�#�2H��T�Br��o��5;��4˸��K�nQ���$�r�u�;���o��؉�w���0���r8	K~\�^����Ly��)n/�g���[K����$w�<�e���Hq�÷L6n�����;�ɻ��M2Ycx�sro��5��F��o�@zt�5�&�����]rD$K~�����뭸��z�o㒙�Q|�dw����ݑa�֒.y0�p+��d83�dkI��mĉ��tWz���̒�%YrO���6^�с�%[K��k\'3���s K�,9����s�}H�1`7v;Sqgɣ1��=�Q��x����d����xDbR%{�J�X��]�XIz?���3Y���`o4&5�$K���V�+�bsk��n5�m�$�㽃�O'���Csr|��d9Y�+!�Q���>��z*$��G����9���'�ة��J{KH��v*�G��CT��g�����PN����n�H�;M����Ãcp����� Ǉ�%v�9��Yi����"��ʸdqFǟi�L89�/B�d��������n�b�H�ٚ��,q�0_�K���;އe�Lq�S$��֙L��H���3���H�Sr�`�9�%� ��Xr���b��wD�m�7�)��Kgߨ`rvA�����ߩd����J�i�_�d�=���
&�;��F����_�v2�:�����{�qk�*nu��FK�<ɯ�WW���F�Yr�G#٭�z�[�K��h$�ō�N�����L׭��ve���-���,Ya��ש[s�����{�JE����%GȪ��(H�Nv���AK��Q�?H_��.=�`�2*9�F�$�I���,�
&,9K��K6`�,9�%,�%G`�T0a�1X2�X�Kf�!,�`�,9K��	K����d��X2Ka�Kf�X2LXr�L%�l��YrK&X2K����`c�d*�d�̒CX2��Yr��H>?K�~��g��X�S��f��3����oI�U�Q��~����O�~�}���5O�!,�`�,9K��	K����d��X2Ka�Kf�X2LXr�L%�l��YrK&X2K����`c�d*�d�̒CX2��Yr�L��%Sɀ%�d�	�̒#�d*���,�J,ـ%��4��(�%Gx��˿�$��˿�k��$��D�;���
�$_'�D��պ�$'�.K��d��%S��%ǰC��$ξQ�$����
&�ߩ`p�V}J%��i�T0��Q���{�N&V��d��D2����s K�,9����s�ϑ�������~%���B�m����-y�@HN���<'G����E�hxp|r��d���.���E�8)|��:S|J���$y8�~:�����pr��w�<���-g������w�X>88:��d��#1W'8��d������Ӈ�C��7Jt|g���ј�
���A2��d��^$3ن%� ��Xr`�9�%� ��Xr`�9��?�c�I���K~���*�qk�#��Aޓ$�֒�bS4;0�Ḇ$�����[&����$�>����d��}M��wC�$�5�����h�&�����d�Xr`�9����yK�a��ϗo���j�d�e�6����ɟI�d�l!i�S%�e�Hu�.�}�=����i�/��d��5y�s��W�x%����^�%<����-#�K$_A�y%+�����Z.�ѿ��K�WңԇĒ���k��ۿ��Kf�aB�W�*�Ks5�b�N���Riv�N�@K���*1͚�^"�ղ֬$�ej_V2�1C
�)�$ɾ�H01���"�Ĭ���=9��q��gl�q,4:�4��R2 ��km��9le��CuN��ץf<�d� �+�ʧe���괤��2D8a�d囲M���M��t`:F�8�Ἃ�a��M �e|cu��U9Xk�%��ejp��������PЂfd����M����m�YwbB���Q2��1��8�"P�>%���p��P G@��c,�ku�$h@<#P2.�ש��|G �,a�����Vp)��qY���r��2�.�5��,@�@=J����t������Z]D��=-��I2�j������m<��D���l
�8T�n���NcU�z���
z�Iț�$9b�[�� �������48�36�͒DAI��Ғŵ����3|��f�s8\������a��}6l?~�n�SlHf',9}�q����;"(��0�    IEND�B`�PK
     ąnY)t8A�  �  /   images/d8a1d1b0-d05e-462a-97fe-7e9bb74087a2.png�PNG

   IHDR  �   �   @w��   gAMA  ���a   �PLTEZs(z4�ǩYYY=H'��3zi���'''Ne$r�,X�O=�O(O0���>>>x��Z�j$7(��i:ZAm�." 000+}:{�1Xa�˸��4�����d@�C*+,j�VRRRb�)I\%f�t����jjj~�1���Th)�`$=*������III���L�Hbbc5�@��lv�.BBB��ivxv��ov�\���)k5s��b�S������osk��e��̴ӻ���o�Y~��������N���   	pHYs  �  ��o�d  �IDATx��[���\;����HYA`FW��p�OW�
:|��sۤI��`CSHl~��M����INNC�;����6�x��oN�f?a]�7'x�-n����~Û��5<PwC�i�Si��},�����x��oV񦛰���	ޜ��#���C�Nܺ�6H�=���ov����������d�ƭ?��A�;��M0R�����:f� �lNa#����W�9~x0���'
�yp��kZc�pC�1d��ŭC��ލ!{�� ?�ݣ�ڍB^X��2�!w7重����ި&�����=�톐���B�/��?!d�7�F�k��޳60dd� ��ֽ�5�lx��?�����Cٷ�m`��A~��v���f�v0䘵�2�^��E�2��v�$񗷷���H`���_;��2��MX����E��5���;q������F��Cv�p7�|T�X�=�����QkZ��B�8Q�F��{�q�����v�b��T�� ��1<�2�8Ɛ��d7�F�ae���{qk#f� ��:�l��}��ŭ'$k7n-�L'�р�!��ƹ:]9���B�'�A>���p�1��ؓ�8�[
� �a��W ��q�2��Ɛ�D�%TU=��>C��C�`��l��9��@�/�� �FprИ�}�MX��kh����A��ؓ�u/n� �G�{���60��A>���no�A�с�(f-���� c�p� d��i#9IW���/�/_"ѵ�r��1��� ��#�s��/���%]{��	k��ŭ;�5
�l� ��F�HZ;q���g�Ñ��G��Y�B�z�0�Ydu��!/�d�#ox����p�	��p` �S�	Ν���٩�ֺO��St���):|��&x���)�z��N�=����! ٍ�l���@�jlb��>�0�Ü s��0���_p*eB��S��a�B�5�����
)b�Ӹ��I)p�g!�: ��q���D����A�A�5�-n��S�5�+�Ԥ�mD1a�A܈�WSY#���@�8T��I)p.��F�T:�X����2@��'��FN��ck�hqFq���EߎY��^o="Y��oG7a��=v�d-)c9���� ����w�F�{4��Tfg;�����ڌ[k	k{�ֲ"��A�q�A.:��t\*��8�b|F��\��}���J��E�&<�~
@�1j0�n��pD�YD�"� �0�-�x�h��,��*t���-8�[�`��*��'=N��pMMI>SDs���*��|a��ZNMcQ�]O�^l��+�$S5�����4dea��D�q�6LE�u�o��T�d��9�M&�j$�J�$WInm�|(�@�0�Oú��=kO���Yk�#m���aj{CM�3{��ꃣ���r���T�����/M{}מ�Ŭ�A~���%����i8�-Jsr������%�t��zO�-��A;�Ɋ�t�R�!�/Jm���p����Q���Z?ռ���b,�(�����XR�|%��D��XVݜ���U�eUz�+�|z�w����=OO��o��^uJ�*AycO.�)	��!wW ��J"�C�iw��ɍc%1UN@�ȓ�j��ɍ������H�]_���^,f}9+�zr���u[ԃ�8.w�t�iZ�m�G���uh�kj�,��ɂdmY���|^\��d%yD�<�/�RI3M��)O�X��Z{jϽ��^<�m[y��"{�Џ�=6�˹Y,�ʓeV�ܵ�,���B}~)O.��������/���1��$�h�2G�ݲ�8"s���⃋����8h�)S!��R�V*�5�V"^O��O.*?�(���J�[N�]�W�J��E����k��K�'�*?�*���e�U�ҠV����P��gO.7*��vKo)�^��A豩��R�݃<����������O��N!E����L���^��O~�-�uʘ\��3n��D���g9��oL.���|Y���'ѓ�8rKI�]��C�?��奭]ִٓ��Z��"�"��r�ސ��Y4��r�d��$��A�y���R� � ��P>c��,�r��d��ٓ
��b�\{����vi�x�nYVs�ӋWK�-b�E+�r+�[��ә���P۾�����c<��j��|��aL��)źE(� 
�����ux؈�dk�l�S��2{��ńBJۛ��=|t�vY<��Z 9�'��z���-J�(��l� 3Sߛ$cz#ӿ��5�5�@�J�!�ԪI����&��"�,J�h�S\�|Zt6�%�"՚Ԙ5m'�����kr�^[^.��wFO����Ei��T����ʞh��������iyY:������|�I����~�~���l�V�ʞCw�g�d"d�5/K��j��Y*��/��ؓ�.�Ij)S�-6��v���HZ����&E��d�M7&�#��ƥ�.\�I.�c(fQ3x�	&�+�Ry�� �.A,f���t׌c2Cq�1��]#Y �g :�Pͥ�;�)�5��j��:�l=[�$zw��1^Y�ə 7X�kݵ��5Kwme�d}g�̥�f�ŉ�Y3^�JHƻ�i�C�8�$�D�D����x29��/w-~t�%)ؘL����=.c�8�5�'g�x�]�8O&��Ǥ�t�ۏ�y���D�9d�䊮E�Ԙ[t-kt-Nw-Btݒ<��sL�*���R�c���y2[w�b���٣kI2^,����]3�,��q�Q�1��PJ�����|�jb��/����r�]�-Mc�ŭ<�$��d�s��J����n�K�a�K��5��]g^㵻1���<9��aBl%�%m'3EןqLfhh�cr�񘊮YZ�gt��'[\2^��䮛,��Eגd��>w�4�b�xmu���]�Y*�>�L<F�s��e��D�b��-�$>��Й�yv�����z�)��O�I�N|����:͜�n��|���&�H�؎�~ܻ�l���D�>���ߌ?�]P���0MB9�OpOB��R�ץ�R��0�:�=]V�[��wчO�J�\ھ��/��kޡ��lƞ|�4��)}�Wr�E]�ƣ�y{r�i� ���Pb�΅�������h�� ��L49�)�,�|����dkƋ<c��<Y�K�l���糷����*�`�L�J���x�x1Y��ӕ�<s�;Hk��ƫ��%��	t�Kt�d(�deH��fmZ��u�\���x1]��se�.>AA~E�Wkv�F�"��j�}�����]L��ş1��n9��u�W��8�5^,)�A�~t��yrnѵՒxL��g�r�BQ��7R��'�"��ݵPw�IomeLf���N�x��	�xQ�dʡs�������͓ڟ�5s�
��R�.��>&S�OP�������]�]K<&�H�#w-otm��ae��%��P<<Y�1�G2����/�*J�T*��d���ԧ��w�ٵ''����U(Q�dѣ�c�/&�'�?>�q=������1��~�1�'�|��I����W��k._H�r���D�Y�Z���M�9���E�-�W&O�|2	r7OfiQ��E�'��Y ��dJ�D�'7Y���,T�5�K��{���Ა�ϧ�ӓ�X�L��<�	��E$kz1�b���� � V�i�Mm$�I��ȍl�ZC,�јL�{��,�:�,{��ۚ�,�Lƌ��<�l�uZO�@�_����brʹ�4�Lu�=>��/�2624؊'�;�6m=��Ӗ�kͳ!^��k+cr1ĥ�y���D����)(�;PW�\ mqLVڑ�]+�D���
�h��zr�|P� [-%�t������F�G��$�~TVg���A��M��$��|#�֙�ɍr���7���p�b�q&O�(�T����}��R{��H�����8�'{������P��Q�k7y*ǪEӏ}R_�ٓ=�哃ʅG��Үuq� 2���?�RFdDY=r�>�j�=x)�:�^4��^��재$��x���R�\ )O.��'@ʓ �����Hyr���˧Jb*���ܓO�����@�<�7��=%au�ɓ�~]JBjo��'����7�����'���E�m����i��c�^�C�7��2����u{�M����'��˓��XèOd����k��#e9�h����n�ʲ�'@*�U )O.��'@�=���MCIF�|%�B�r�ܯʗe�ͿD����+_�P�T�ʗ��1��,����@�nH���#���Huk��E�m�w0�j�SI��|�k���=��K ]'4^��0�k~�?<�?�$�@�@�v{�^�s��^v�C}����=�PCm���0�<ss�J�(���n�mdjJ2ˮN��ɴ�`��Ը4U��U��0�3�l���[S�S���^P@����[��)ɨ^���B�&�c�qH�P=��
����#/(�����Z���G��MS�N&D<�gկ3xd0>C�n�U�J�W�Y��
w� 2��G�Zy]I&�K�q\�wd?�v"	4��]MI2u��.��#-��C��@��)I������� �m�#�s%�F��%'�+�	��$� �e���d�0&��d��<�8�Z �ޯx�F�,Q�G`�q�+4�;��ʔ��6�0��~9�x���� �����Jr	��h�l��:�܁	���+��V�,��eF����f5a�#�
5�_��������109��'O�Ϡز |���W����$��Iȸ��Y�5^Uأ�U��Y�7�o��jM��؊���;�ؕb�$� R���y]���8��#�[    IEND�B`�PK 
     ąnY�|oy[ y[                  cirkitFile.jsonPK 
     ąnY                        �[ jsons/PK 
     ąnYc�E�  �               �[ jsons/user_defined.jsonPK 
     ąnY                        �u images/PK 
     ąnY�m�ځ ځ /             "v images/1c49e1bc-8662-4f8f-9dd9-28b8f22266b8.pngPK 
     ąnY���T0  T0  /             I� images/5107842f-df24-4ed4-8dc8-476b8a0f3ddf.pngPK 
     ąnYP��/ǽ  ǽ  /             �( images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     ąnY$7h�!  �!  /             �� images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     ąnY��ƌ  �  /             <	 images/04d2d11f-9dbd-4a2c-b6c9-835d97151b37.pngPK 
     ąnY)t8A�  �  /              images/d8a1d1b0-d05e-462a-97fe-7e9bb74087a2.pngPK    
 
   :.   